.SUBCKT MULTIPLIER_G4_12_7685 A B C Y VCC GND
Mcl0ECICH_0#0 cl0ECICH_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_0#1 cl0ECICH_0#Y C GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#0 VCC B cl0ECICH_1#clCZWK1K_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#1 cl0ECICH_1#clCZWK1K_0#a_18_54# cl0ECICH_1#clCZWK1K_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#2 cl0ECICH_1#clCZWK1K_0#Y cl0ECICH_1#clCZWK1K_0#a_2_6# cl0ECICH_1#clCZWK1K_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#3 cl0ECICH_1#clCZWK1K_0#a_35_54# B cl0ECICH_1#clCZWK1K_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#4 VCC A cl0ECICH_1#clCZWK1K_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#5 cl0ECICH_1#clCZWK1K_0#a_12_41# A VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#6 GND B cl0ECICH_1#clCZWK1K_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#7 cl0ECICH_1#clCZWK1K_0#a_18_6# cl0ECICH_1#clCZWK1K_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#8 cl0ECICH_1#clCZWK1K_0#Y B cl0ECICH_1#clCZWK1K_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#9 cl0ECICH_1#clCZWK1K_0#a_35_6# cl0ECICH_1#clCZWK1K_0#a_2_6# cl0ECICH_1#clCZWK1K_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#10 GND A cl0ECICH_1#clCZWK1K_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_0#11 cl0ECICH_1#clCZWK1K_0#a_12_41# A GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#0 VCC cl0ECICH_1#clCZWK1K_0#Y cl0ECICH_1#clCZWK1K_1#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#1 cl0ECICH_1#clCZWK1K_1#a_18_54# cl0ECICH_1#clCZWK1K_1#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#2 Y cl0ECICH_1#clCZWK1K_1#a_2_6# cl0ECICH_1#clCZWK1K_1#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#3 cl0ECICH_1#clCZWK1K_1#a_35_54# cl0ECICH_1#clCZWK1K_0#Y Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#4 VCC cl0ECICH_0#Y cl0ECICH_1#clCZWK1K_1#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#5 cl0ECICH_1#clCZWK1K_1#a_12_41# cl0ECICH_0#Y VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#6 GND cl0ECICH_1#clCZWK1K_0#Y cl0ECICH_1#clCZWK1K_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#7 cl0ECICH_1#clCZWK1K_1#a_18_6# cl0ECICH_1#clCZWK1K_1#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#8 Y cl0ECICH_1#clCZWK1K_0#Y cl0ECICH_1#clCZWK1K_1#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#9 cl0ECICH_1#clCZWK1K_1#a_35_6# cl0ECICH_1#clCZWK1K_1#a_2_6# Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#10 GND cl0ECICH_0#Y cl0ECICH_1#clCZWK1K_1#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0ECICH_1#clCZWK1K_1#11 cl0ECICH_1#clCZWK1K_1#a_12_41# cl0ECICH_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 3|3|MULTIPLIER_G1_25_27|INVX1=1|INPUT:Y-INVX1:A=1|INPUT:Y-MULTIPLIER_G1_25_27:A,B,C=2|INVX1:Y-MULTIPLIER_G1_25_27:A,B,C=1|11110
* 538 occurrences in design
* each contains 2 cells
* pin map: {'n7847': 'A', 'n7842': 'B', 'x2': 'C'} {'n7848': 'Y'}
* function: (A&B&~C)|(A&C&~B)|(B&C&~A)|(~A&~B&~C)
* Example occurence:
*   .subckt INVX1 A=x2 Y=n132
*   .subckt MULTIPLIER_G1_25_27 A=n132 B=n7842 C=n7847 Y=n7848
