.SUBCKT BAR_G3_4_5 A B C VDD VSS Y
Mcl2ZSDQD_0#M0 cl2ZSDQD_0#Y C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_0#M1 cl2ZSDQD_0#Y C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_1#clJZI4Y2_0#M3 cl2ZSDQD_1#clJZI4Y2_0#net16 A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
Mcl2ZSDQD_1#clJZI4Y2_0#M2 cl2ZSDQD_1#clJZI4Y2_0#Y B cl2ZSDQD_1#clJZI4Y2_0#net16 VSS nmos_lvt w=162.00n l=20n nfin=6
Mcl2ZSDQD_1#clJZI4Y2_0#M1 cl2ZSDQD_1#clJZI4Y2_0#Y B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_1#clJZI4Y2_0#M0 cl2ZSDQD_1#clJZI4Y2_0#Y A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#M5 VSS cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net7 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#Y VSS nmos_lvt w=162.00n l=20n nfin=6
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#M1 VSS cl2ZSDQD_1#clJZI4Y2_1#C cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net7 VSS nmos_lvt w=54.0n l=20n nfin=2
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#M2 VSS cl2ZSDQD_0#Y cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net7 VSS nmos_lvt w=54.0n l=20n nfin=2
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#M0 VDD cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net7 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#Y VDD pmos_lvt w=162.00n l=20n nfin=6
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#M4 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net15 cl2ZSDQD_1#clJZI4Y2_1#C cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net7 VDD pmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#M3 VDD cl2ZSDQD_0#Y cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#net15 VDD pmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#M4 Y cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net10 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#M1 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net10 cl2ZSDQD_1#clJZI4Y2_0#Y VDD VDD pmos_lvt w=54.0n l=20n nfin=2
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#M0 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net10 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#Y VDD VDD pmos_lvt w=54.0n l=20n nfin=2
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#M5 Y cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net10 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#M3 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net20 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_0#Y VSS VSS nmos_lvt w=81.0n l=20n nfin=3
Mcl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#M2 cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net10 cl2ZSDQD_1#clJZI4Y2_0#Y cl2ZSDQD_1#clJZI4Y2_1#clTAMZRU_1#net20 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS 
* pattern code: 4|3|BAR_G2_3_5|INVx1=1|INPUT:Y-BAR_G2_3_5:B=1|INPUT:Y-BAR_G2_3_5:C=1|INPUT:Y-INVx1:A=1|INVx1:Y-BAR_G2_3_5:A=1|01111
* 96 occurrences in design
* each contains 2 cells
* function: (B&~A)|(~B&~C)
* Example occurence:
*   .subckt INVx1 A=x60 Y=n190
*   .subckt BAR_G2_3_5 A=n190 B=x128 C=x59 Y=n359
