.SUBCKT MULTIPLIER_G3_77_78 A B C D Y VCC GND
Mcl7XSHR2_0#0 VCC C cl7XSHR2_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#1 cl7XSHR2_0#a_18_54# cl7XSHR2_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#2 cl7XSHR2_0#Y cl7XSHR2_0#a_2_6# cl7XSHR2_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#3 cl7XSHR2_0#a_35_54# C cl7XSHR2_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#4 VCC D cl7XSHR2_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#5 cl7XSHR2_0#a_12_41# D VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#6 GND C cl7XSHR2_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#7 cl7XSHR2_0#a_18_6# cl7XSHR2_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#8 cl7XSHR2_0#Y C cl7XSHR2_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#9 cl7XSHR2_0#a_35_6# cl7XSHR2_0#a_2_6# cl7XSHR2_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#10 GND D cl7XSHR2_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_0#11 cl7XSHR2_0#a_12_41# D GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#0 VCC A cl7XSHR2_1#clCZWK1K_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#1 cl7XSHR2_1#clCZWK1K_0#a_18_54# cl7XSHR2_1#clCZWK1K_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#2 cl7XSHR2_1#clCZWK1K_0#Y cl7XSHR2_1#clCZWK1K_0#a_2_6# cl7XSHR2_1#clCZWK1K_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#3 cl7XSHR2_1#clCZWK1K_0#a_35_54# A cl7XSHR2_1#clCZWK1K_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#4 VCC cl7XSHR2_0#Y cl7XSHR2_1#clCZWK1K_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#5 cl7XSHR2_1#clCZWK1K_0#a_12_41# cl7XSHR2_0#Y VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#6 GND A cl7XSHR2_1#clCZWK1K_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#7 cl7XSHR2_1#clCZWK1K_0#a_18_6# cl7XSHR2_1#clCZWK1K_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#8 cl7XSHR2_1#clCZWK1K_0#Y A cl7XSHR2_1#clCZWK1K_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#9 cl7XSHR2_1#clCZWK1K_0#a_35_6# cl7XSHR2_1#clCZWK1K_0#a_2_6# cl7XSHR2_1#clCZWK1K_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#10 GND cl7XSHR2_0#Y cl7XSHR2_1#clCZWK1K_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_0#11 cl7XSHR2_1#clCZWK1K_0#a_12_41# cl7XSHR2_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#0 VCC cl7XSHR2_1#clCZWK1K_0#Y cl7XSHR2_1#clCZWK1K_1#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#1 cl7XSHR2_1#clCZWK1K_1#a_18_54# cl7XSHR2_1#clCZWK1K_1#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#2 Y cl7XSHR2_1#clCZWK1K_1#a_2_6# cl7XSHR2_1#clCZWK1K_1#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#3 cl7XSHR2_1#clCZWK1K_1#a_35_54# cl7XSHR2_1#clCZWK1K_0#Y Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#4 VCC B cl7XSHR2_1#clCZWK1K_1#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#5 cl7XSHR2_1#clCZWK1K_1#a_12_41# B VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#6 GND cl7XSHR2_1#clCZWK1K_0#Y cl7XSHR2_1#clCZWK1K_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#7 cl7XSHR2_1#clCZWK1K_1#a_18_6# cl7XSHR2_1#clCZWK1K_1#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#8 Y cl7XSHR2_1#clCZWK1K_0#Y cl7XSHR2_1#clCZWK1K_1#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#9 cl7XSHR2_1#clCZWK1K_1#a_35_6# cl7XSHR2_1#clCZWK1K_1#a_2_6# Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#10 GND B cl7XSHR2_1#clCZWK1K_1#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl7XSHR2_1#clCZWK1K_1#11 cl7XSHR2_1#clCZWK1K_1#a_12_41# B GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 3|4|MULTIPLIER_G1_25_27|XNOR2X1=1|INPUT:Y-MULTIPLIER_G1_25_27:A,B,C=2|INPUT:Y-XNOR2X1:A,B=2|XNOR2X1:Y-MULTIPLIER_G1_25_27:A,B,C=1|111101
* 1020 occurrences in design
* each contains 2 cells
* pin map: {'n330': 'A', 'n333': 'B', 'n132': 'C', 'n313': 'D'} {'y4': 'Y'}
* function: (A&B&C&D)|(A&B&~C&~D)|(A&C&~B&~D)|(A&D&~B&~C)|(B&C&~A&~D)|(B&D&~A&~C)|(C&D&~A&~B)|(~A&~B&~C&~D)
* Example occurence:
*   .subckt XNOR2X1 A=n132 B=n313 Y=n314
*   .subckt MULTIPLIER_G1_25_27 A=n333 B=n330 C=n314 Y=y4
