.SUBCKT CTRL_G1_68_69 A B C Y VCC GND
Mcl0E90G9_0#0 cl0E90G9_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_0#1 VCC A cl0E90G9_0#Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_0#2 cl0E90G9_0#Y B VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_0#3 cl0E90G9_0#a_9_6# C GND GND nmos w=0.75u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_0#4 cl0E90G9_0#a_14_6# A cl0E90G9_0#a_9_6# GND nmos w=0.75u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_0#5 cl0E90G9_0#Y B cl0E90G9_0#a_14_6# GND nmos w=0.75u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_1#0 Y cl0E90G9_0#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0E90G9_1#1 Y cl0E90G9_0#Y GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 2|3|INVX1|NAND3X1=1|INPUT:Y-NAND3X1:A,B,C=3|NAND3X1:Y-INVX1:A=1|11101
* 4 occurrences in design
* each contains 2 cells
* pin map: {'n10': 'A', 'n76': 'B', 'n9': 'C'} {'y11': 'Y'}
* function: A&B&C
* Example occurence:
*   .subckt NAND3X1 A=n9 B=n10 C=n76 Y=n77
*   .subckt INVX1 A=n77 Y=y11
