// Benchmark "benchmark/aig/full_adder_256" written by ABC on Tue Jan  2 21:13:28 2024

module ADDER_G0_20_21  ( A, B, C, Y );
  input A,B,C;
  output Y;
  assign Y=(A*B*C)+(A*!B*!C)+(B*!A*!C)+(C*!A*!B);
endmodule

module ADDER_G2_27_28_29  ( A, B, C, Y );
  input A,B,C;
  output Y;
  assign Y=(A*B)+(A*C)+(B*C);
endmodule

module full_adder_256  ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511, pi512,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511, pi512;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256;
  wire new_n772_, new_n774_, new_n776_, new_n778_, new_n780_, new_n782_,
    new_n784_, new_n786_, new_n788_, new_n790_, new_n792_, new_n794_,
    new_n796_, new_n798_, new_n800_, new_n802_, new_n804_, new_n806_,
    new_n808_, new_n810_, new_n812_, new_n814_, new_n816_, new_n818_,
    new_n820_, new_n822_, new_n824_, new_n826_, new_n828_, new_n830_,
    new_n832_, new_n834_, new_n836_, new_n838_, new_n840_, new_n842_,
    new_n844_, new_n846_, new_n848_, new_n850_, new_n852_, new_n854_,
    new_n856_, new_n858_, new_n860_, new_n862_, new_n864_, new_n866_,
    new_n868_, new_n870_, new_n872_, new_n874_, new_n876_, new_n878_,
    new_n880_, new_n882_, new_n884_, new_n886_, new_n888_, new_n890_,
    new_n892_, new_n894_, new_n896_, new_n898_, new_n900_, new_n902_,
    new_n904_, new_n906_, new_n908_, new_n910_, new_n912_, new_n914_,
    new_n916_, new_n918_, new_n920_, new_n922_, new_n924_, new_n926_,
    new_n928_, new_n930_, new_n932_, new_n934_, new_n936_, new_n938_,
    new_n940_, new_n942_, new_n944_, new_n946_, new_n948_, new_n950_,
    new_n952_, new_n954_, new_n956_, new_n958_, new_n960_, new_n962_,
    new_n964_, new_n966_, new_n968_, new_n970_, new_n972_, new_n974_,
    new_n976_, new_n978_, new_n980_, new_n982_, new_n984_, new_n986_,
    new_n988_, new_n990_, new_n992_, new_n994_, new_n996_, new_n998_,
    new_n1000_, new_n1002_, new_n1004_, new_n1006_, new_n1008_, new_n1010_,
    new_n1012_, new_n1014_, new_n1016_, new_n1018_, new_n1020_, new_n1022_,
    new_n1024_, new_n1026_, new_n1028_, new_n1030_, new_n1032_, new_n1034_,
    new_n1036_, new_n1038_, new_n1040_, new_n1042_, new_n1044_, new_n1046_,
    new_n1048_, new_n1050_, new_n1052_, new_n1054_, new_n1056_, new_n1058_,
    new_n1060_, new_n1062_, new_n1064_, new_n1066_, new_n1068_, new_n1070_,
    new_n1072_, new_n1074_, new_n1076_, new_n1078_, new_n1080_, new_n1082_,
    new_n1084_, new_n1086_, new_n1088_, new_n1090_, new_n1092_, new_n1094_,
    new_n1096_, new_n1098_, new_n1100_, new_n1102_, new_n1104_, new_n1106_,
    new_n1108_, new_n1110_, new_n1112_, new_n1114_, new_n1116_, new_n1118_,
    new_n1120_, new_n1122_, new_n1124_, new_n1126_, new_n1128_, new_n1130_,
    new_n1132_, new_n1134_, new_n1136_, new_n1138_, new_n1140_, new_n1142_,
    new_n1144_, new_n1146_, new_n1148_, new_n1150_, new_n1152_, new_n1154_,
    new_n1156_, new_n1158_, new_n1160_, new_n1162_, new_n1164_, new_n1166_,
    new_n1168_, new_n1170_, new_n1172_, new_n1174_, new_n1176_, new_n1178_,
    new_n1180_, new_n1182_, new_n1184_, new_n1186_, new_n1188_, new_n1190_,
    new_n1192_, new_n1194_, new_n1196_, new_n1198_, new_n1200_, new_n1202_,
    new_n1204_, new_n1206_, new_n1208_, new_n1210_, new_n1212_, new_n1214_,
    new_n1216_, new_n1218_, new_n1220_, new_n1222_, new_n1224_, new_n1226_,
    new_n1228_, new_n1230_, new_n1232_, new_n1234_, new_n1236_, new_n1238_,
    new_n1240_, new_n1242_, new_n1244_, new_n1246_, new_n1248_, new_n1250_,
    new_n1252_, new_n1254_, new_n1256_, new_n1258_, new_n1260_, new_n1262_,
    new_n1264_, new_n1266_, new_n1268_, new_n1270_, new_n1272_, new_n1274_,
    new_n1276_, new_n1278_, new_n1280_;
  ADDER_G0_20_21    g000(.A(pi512), .B(pi256), .C(pi000), .Y(po000));
  ADDER_G2_27_28_29 g001(.A(pi512), .B(pi256), .C(pi000), .Y(new_n772_));
  ADDER_G0_20_21    g002(.A(new_n772_), .B(pi257), .C(pi001), .Y(po001));
  ADDER_G2_27_28_29 g003(.A(new_n772_), .B(pi257), .C(pi001), .Y(new_n774_));
  ADDER_G0_20_21    g004(.A(new_n774_), .B(pi258), .C(pi002), .Y(po002));
  ADDER_G2_27_28_29 g005(.A(new_n774_), .B(pi258), .C(pi002), .Y(new_n776_));
  ADDER_G0_20_21    g006(.A(new_n776_), .B(pi259), .C(pi003), .Y(po003));
  ADDER_G2_27_28_29 g007(.A(new_n776_), .B(pi259), .C(pi003), .Y(new_n778_));
  ADDER_G0_20_21    g008(.A(new_n778_), .B(pi260), .C(pi004), .Y(po004));
  ADDER_G2_27_28_29 g009(.A(new_n778_), .B(pi260), .C(pi004), .Y(new_n780_));
  ADDER_G0_20_21    g010(.A(new_n780_), .B(pi261), .C(pi005), .Y(po005));
  ADDER_G2_27_28_29 g011(.A(new_n780_), .B(pi261), .C(pi005), .Y(new_n782_));
  ADDER_G0_20_21    g012(.A(new_n782_), .B(pi262), .C(pi006), .Y(po006));
  ADDER_G2_27_28_29 g013(.A(new_n782_), .B(pi262), .C(pi006), .Y(new_n784_));
  ADDER_G0_20_21    g014(.A(new_n784_), .B(pi263), .C(pi007), .Y(po007));
  ADDER_G2_27_28_29 g015(.A(new_n784_), .B(pi263), .C(pi007), .Y(new_n786_));
  ADDER_G0_20_21    g016(.A(new_n786_), .B(pi264), .C(pi008), .Y(po008));
  ADDER_G2_27_28_29 g017(.A(new_n786_), .B(pi264), .C(pi008), .Y(new_n788_));
  ADDER_G0_20_21    g018(.A(new_n788_), .B(pi265), .C(pi009), .Y(po009));
  ADDER_G2_27_28_29 g019(.A(new_n788_), .B(pi265), .C(pi009), .Y(new_n790_));
  ADDER_G0_20_21    g020(.A(new_n790_), .B(pi266), .C(pi010), .Y(po010));
  ADDER_G2_27_28_29 g021(.A(new_n790_), .B(pi266), .C(pi010), .Y(new_n792_));
  ADDER_G0_20_21    g022(.A(new_n792_), .B(pi267), .C(pi011), .Y(po011));
  ADDER_G2_27_28_29 g023(.A(new_n792_), .B(pi267), .C(pi011), .Y(new_n794_));
  ADDER_G0_20_21    g024(.A(new_n794_), .B(pi268), .C(pi012), .Y(po012));
  ADDER_G2_27_28_29 g025(.A(new_n794_), .B(pi268), .C(pi012), .Y(new_n796_));
  ADDER_G0_20_21    g026(.A(new_n796_), .B(pi269), .C(pi013), .Y(po013));
  ADDER_G2_27_28_29 g027(.A(new_n796_), .B(pi269), .C(pi013), .Y(new_n798_));
  ADDER_G0_20_21    g028(.A(new_n798_), .B(pi270), .C(pi014), .Y(po014));
  ADDER_G2_27_28_29 g029(.A(new_n798_), .B(pi270), .C(pi014), .Y(new_n800_));
  ADDER_G0_20_21    g030(.A(new_n800_), .B(pi271), .C(pi015), .Y(po015));
  ADDER_G2_27_28_29 g031(.A(new_n800_), .B(pi271), .C(pi015), .Y(new_n802_));
  ADDER_G0_20_21    g032(.A(new_n802_), .B(pi272), .C(pi016), .Y(po016));
  ADDER_G2_27_28_29 g033(.A(new_n802_), .B(pi272), .C(pi016), .Y(new_n804_));
  ADDER_G0_20_21    g034(.A(new_n804_), .B(pi273), .C(pi017), .Y(po017));
  ADDER_G2_27_28_29 g035(.A(new_n804_), .B(pi273), .C(pi017), .Y(new_n806_));
  ADDER_G0_20_21    g036(.A(new_n806_), .B(pi274), .C(pi018), .Y(po018));
  ADDER_G2_27_28_29 g037(.A(new_n806_), .B(pi274), .C(pi018), .Y(new_n808_));
  ADDER_G0_20_21    g038(.A(new_n808_), .B(pi275), .C(pi019), .Y(po019));
  ADDER_G2_27_28_29 g039(.A(new_n808_), .B(pi275), .C(pi019), .Y(new_n810_));
  ADDER_G0_20_21    g040(.A(new_n810_), .B(pi276), .C(pi020), .Y(po020));
  ADDER_G2_27_28_29 g041(.A(new_n810_), .B(pi276), .C(pi020), .Y(new_n812_));
  ADDER_G0_20_21    g042(.A(new_n812_), .B(pi277), .C(pi021), .Y(po021));
  ADDER_G2_27_28_29 g043(.A(new_n812_), .B(pi277), .C(pi021), .Y(new_n814_));
  ADDER_G0_20_21    g044(.A(new_n814_), .B(pi278), .C(pi022), .Y(po022));
  ADDER_G2_27_28_29 g045(.A(new_n814_), .B(pi278), .C(pi022), .Y(new_n816_));
  ADDER_G0_20_21    g046(.A(new_n816_), .B(pi279), .C(pi023), .Y(po023));
  ADDER_G2_27_28_29 g047(.A(new_n816_), .B(pi279), .C(pi023), .Y(new_n818_));
  ADDER_G0_20_21    g048(.A(new_n818_), .B(pi280), .C(pi024), .Y(po024));
  ADDER_G2_27_28_29 g049(.A(new_n818_), .B(pi280), .C(pi024), .Y(new_n820_));
  ADDER_G0_20_21    g050(.A(new_n820_), .B(pi281), .C(pi025), .Y(po025));
  ADDER_G2_27_28_29 g051(.A(new_n820_), .B(pi281), .C(pi025), .Y(new_n822_));
  ADDER_G0_20_21    g052(.A(new_n822_), .B(pi282), .C(pi026), .Y(po026));
  ADDER_G2_27_28_29 g053(.A(new_n822_), .B(pi282), .C(pi026), .Y(new_n824_));
  ADDER_G0_20_21    g054(.A(new_n824_), .B(pi283), .C(pi027), .Y(po027));
  ADDER_G2_27_28_29 g055(.A(new_n824_), .B(pi283), .C(pi027), .Y(new_n826_));
  ADDER_G0_20_21    g056(.A(new_n826_), .B(pi284), .C(pi028), .Y(po028));
  ADDER_G2_27_28_29 g057(.A(new_n826_), .B(pi284), .C(pi028), .Y(new_n828_));
  ADDER_G0_20_21    g058(.A(new_n828_), .B(pi285), .C(pi029), .Y(po029));
  ADDER_G2_27_28_29 g059(.A(new_n828_), .B(pi285), .C(pi029), .Y(new_n830_));
  ADDER_G0_20_21    g060(.A(new_n830_), .B(pi286), .C(pi030), .Y(po030));
  ADDER_G2_27_28_29 g061(.A(new_n830_), .B(pi286), .C(pi030), .Y(new_n832_));
  ADDER_G0_20_21    g062(.A(new_n832_), .B(pi287), .C(pi031), .Y(po031));
  ADDER_G2_27_28_29 g063(.A(new_n832_), .B(pi287), .C(pi031), .Y(new_n834_));
  ADDER_G0_20_21    g064(.A(new_n834_), .B(pi288), .C(pi032), .Y(po032));
  ADDER_G2_27_28_29 g065(.A(new_n834_), .B(pi288), .C(pi032), .Y(new_n836_));
  ADDER_G0_20_21    g066(.A(new_n836_), .B(pi289), .C(pi033), .Y(po033));
  ADDER_G2_27_28_29 g067(.A(new_n836_), .B(pi289), .C(pi033), .Y(new_n838_));
  ADDER_G0_20_21    g068(.A(new_n838_), .B(pi290), .C(pi034), .Y(po034));
  ADDER_G2_27_28_29 g069(.A(new_n838_), .B(pi290), .C(pi034), .Y(new_n840_));
  ADDER_G0_20_21    g070(.A(new_n840_), .B(pi291), .C(pi035), .Y(po035));
  ADDER_G2_27_28_29 g071(.A(new_n840_), .B(pi291), .C(pi035), .Y(new_n842_));
  ADDER_G0_20_21    g072(.A(new_n842_), .B(pi292), .C(pi036), .Y(po036));
  ADDER_G2_27_28_29 g073(.A(new_n842_), .B(pi292), .C(pi036), .Y(new_n844_));
  ADDER_G0_20_21    g074(.A(new_n844_), .B(pi293), .C(pi037), .Y(po037));
  ADDER_G2_27_28_29 g075(.A(new_n844_), .B(pi293), .C(pi037), .Y(new_n846_));
  ADDER_G0_20_21    g076(.A(new_n846_), .B(pi294), .C(pi038), .Y(po038));
  ADDER_G2_27_28_29 g077(.A(new_n846_), .B(pi294), .C(pi038), .Y(new_n848_));
  ADDER_G0_20_21    g078(.A(new_n848_), .B(pi295), .C(pi039), .Y(po039));
  ADDER_G2_27_28_29 g079(.A(new_n848_), .B(pi295), .C(pi039), .Y(new_n850_));
  ADDER_G0_20_21    g080(.A(new_n850_), .B(pi296), .C(pi040), .Y(po040));
  ADDER_G2_27_28_29 g081(.A(new_n850_), .B(pi296), .C(pi040), .Y(new_n852_));
  ADDER_G0_20_21    g082(.A(new_n852_), .B(pi297), .C(pi041), .Y(po041));
  ADDER_G2_27_28_29 g083(.A(new_n852_), .B(pi297), .C(pi041), .Y(new_n854_));
  ADDER_G0_20_21    g084(.A(new_n854_), .B(pi298), .C(pi042), .Y(po042));
  ADDER_G2_27_28_29 g085(.A(new_n854_), .B(pi298), .C(pi042), .Y(new_n856_));
  ADDER_G0_20_21    g086(.A(new_n856_), .B(pi299), .C(pi043), .Y(po043));
  ADDER_G2_27_28_29 g087(.A(new_n856_), .B(pi299), .C(pi043), .Y(new_n858_));
  ADDER_G0_20_21    g088(.A(new_n858_), .B(pi300), .C(pi044), .Y(po044));
  ADDER_G2_27_28_29 g089(.A(new_n858_), .B(pi300), .C(pi044), .Y(new_n860_));
  ADDER_G0_20_21    g090(.A(new_n860_), .B(pi301), .C(pi045), .Y(po045));
  ADDER_G2_27_28_29 g091(.A(new_n860_), .B(pi301), .C(pi045), .Y(new_n862_));
  ADDER_G0_20_21    g092(.A(new_n862_), .B(pi302), .C(pi046), .Y(po046));
  ADDER_G2_27_28_29 g093(.A(new_n862_), .B(pi302), .C(pi046), .Y(new_n864_));
  ADDER_G0_20_21    g094(.A(new_n864_), .B(pi303), .C(pi047), .Y(po047));
  ADDER_G2_27_28_29 g095(.A(new_n864_), .B(pi303), .C(pi047), .Y(new_n866_));
  ADDER_G0_20_21    g096(.A(new_n866_), .B(pi304), .C(pi048), .Y(po048));
  ADDER_G2_27_28_29 g097(.A(new_n866_), .B(pi304), .C(pi048), .Y(new_n868_));
  ADDER_G0_20_21    g098(.A(new_n868_), .B(pi305), .C(pi049), .Y(po049));
  ADDER_G2_27_28_29 g099(.A(new_n868_), .B(pi305), .C(pi049), .Y(new_n870_));
  ADDER_G0_20_21    g100(.A(new_n870_), .B(pi306), .C(pi050), .Y(po050));
  ADDER_G2_27_28_29 g101(.A(new_n870_), .B(pi306), .C(pi050), .Y(new_n872_));
  ADDER_G0_20_21    g102(.A(new_n872_), .B(pi307), .C(pi051), .Y(po051));
  ADDER_G2_27_28_29 g103(.A(new_n872_), .B(pi307), .C(pi051), .Y(new_n874_));
  ADDER_G0_20_21    g104(.A(new_n874_), .B(pi308), .C(pi052), .Y(po052));
  ADDER_G2_27_28_29 g105(.A(new_n874_), .B(pi308), .C(pi052), .Y(new_n876_));
  ADDER_G0_20_21    g106(.A(new_n876_), .B(pi309), .C(pi053), .Y(po053));
  ADDER_G2_27_28_29 g107(.A(new_n876_), .B(pi309), .C(pi053), .Y(new_n878_));
  ADDER_G0_20_21    g108(.A(new_n878_), .B(pi310), .C(pi054), .Y(po054));
  ADDER_G2_27_28_29 g109(.A(new_n878_), .B(pi310), .C(pi054), .Y(new_n880_));
  ADDER_G0_20_21    g110(.A(new_n880_), .B(pi311), .C(pi055), .Y(po055));
  ADDER_G2_27_28_29 g111(.A(new_n880_), .B(pi311), .C(pi055), .Y(new_n882_));
  ADDER_G0_20_21    g112(.A(new_n882_), .B(pi312), .C(pi056), .Y(po056));
  ADDER_G2_27_28_29 g113(.A(new_n882_), .B(pi312), .C(pi056), .Y(new_n884_));
  ADDER_G0_20_21    g114(.A(new_n884_), .B(pi313), .C(pi057), .Y(po057));
  ADDER_G2_27_28_29 g115(.A(new_n884_), .B(pi313), .C(pi057), .Y(new_n886_));
  ADDER_G0_20_21    g116(.A(new_n886_), .B(pi314), .C(pi058), .Y(po058));
  ADDER_G2_27_28_29 g117(.A(new_n886_), .B(pi314), .C(pi058), .Y(new_n888_));
  ADDER_G0_20_21    g118(.A(new_n888_), .B(pi315), .C(pi059), .Y(po059));
  ADDER_G2_27_28_29 g119(.A(new_n888_), .B(pi315), .C(pi059), .Y(new_n890_));
  ADDER_G0_20_21    g120(.A(new_n890_), .B(pi316), .C(pi060), .Y(po060));
  ADDER_G2_27_28_29 g121(.A(new_n890_), .B(pi316), .C(pi060), .Y(new_n892_));
  ADDER_G0_20_21    g122(.A(new_n892_), .B(pi317), .C(pi061), .Y(po061));
  ADDER_G2_27_28_29 g123(.A(new_n892_), .B(pi317), .C(pi061), .Y(new_n894_));
  ADDER_G0_20_21    g124(.A(new_n894_), .B(pi318), .C(pi062), .Y(po062));
  ADDER_G2_27_28_29 g125(.A(new_n894_), .B(pi318), .C(pi062), .Y(new_n896_));
  ADDER_G0_20_21    g126(.A(new_n896_), .B(pi319), .C(pi063), .Y(po063));
  ADDER_G2_27_28_29 g127(.A(new_n896_), .B(pi319), .C(pi063), .Y(new_n898_));
  ADDER_G0_20_21    g128(.A(new_n898_), .B(pi320), .C(pi064), .Y(po064));
  ADDER_G2_27_28_29 g129(.A(new_n898_), .B(pi320), .C(pi064), .Y(new_n900_));
  ADDER_G0_20_21    g130(.A(new_n900_), .B(pi321), .C(pi065), .Y(po065));
  ADDER_G2_27_28_29 g131(.A(new_n900_), .B(pi321), .C(pi065), .Y(new_n902_));
  ADDER_G0_20_21    g132(.A(new_n902_), .B(pi322), .C(pi066), .Y(po066));
  ADDER_G2_27_28_29 g133(.A(new_n902_), .B(pi322), .C(pi066), .Y(new_n904_));
  ADDER_G0_20_21    g134(.A(new_n904_), .B(pi323), .C(pi067), .Y(po067));
  ADDER_G2_27_28_29 g135(.A(new_n904_), .B(pi323), .C(pi067), .Y(new_n906_));
  ADDER_G0_20_21    g136(.A(new_n906_), .B(pi324), .C(pi068), .Y(po068));
  ADDER_G2_27_28_29 g137(.A(new_n906_), .B(pi324), .C(pi068), .Y(new_n908_));
  ADDER_G0_20_21    g138(.A(new_n908_), .B(pi325), .C(pi069), .Y(po069));
  ADDER_G2_27_28_29 g139(.A(new_n908_), .B(pi325), .C(pi069), .Y(new_n910_));
  ADDER_G0_20_21    g140(.A(new_n910_), .B(pi326), .C(pi070), .Y(po070));
  ADDER_G2_27_28_29 g141(.A(new_n910_), .B(pi326), .C(pi070), .Y(new_n912_));
  ADDER_G0_20_21    g142(.A(new_n912_), .B(pi327), .C(pi071), .Y(po071));
  ADDER_G2_27_28_29 g143(.A(new_n912_), .B(pi327), .C(pi071), .Y(new_n914_));
  ADDER_G0_20_21    g144(.A(new_n914_), .B(pi328), .C(pi072), .Y(po072));
  ADDER_G2_27_28_29 g145(.A(new_n914_), .B(pi328), .C(pi072), .Y(new_n916_));
  ADDER_G0_20_21    g146(.A(new_n916_), .B(pi329), .C(pi073), .Y(po073));
  ADDER_G2_27_28_29 g147(.A(new_n916_), .B(pi329), .C(pi073), .Y(new_n918_));
  ADDER_G0_20_21    g148(.A(new_n918_), .B(pi330), .C(pi074), .Y(po074));
  ADDER_G2_27_28_29 g149(.A(new_n918_), .B(pi330), .C(pi074), .Y(new_n920_));
  ADDER_G0_20_21    g150(.A(new_n920_), .B(pi331), .C(pi075), .Y(po075));
  ADDER_G2_27_28_29 g151(.A(new_n920_), .B(pi331), .C(pi075), .Y(new_n922_));
  ADDER_G0_20_21    g152(.A(new_n922_), .B(pi332), .C(pi076), .Y(po076));
  ADDER_G2_27_28_29 g153(.A(new_n922_), .B(pi332), .C(pi076), .Y(new_n924_));
  ADDER_G0_20_21    g154(.A(new_n924_), .B(pi333), .C(pi077), .Y(po077));
  ADDER_G2_27_28_29 g155(.A(new_n924_), .B(pi333), .C(pi077), .Y(new_n926_));
  ADDER_G0_20_21    g156(.A(new_n926_), .B(pi334), .C(pi078), .Y(po078));
  ADDER_G2_27_28_29 g157(.A(new_n926_), .B(pi334), .C(pi078), .Y(new_n928_));
  ADDER_G0_20_21    g158(.A(new_n928_), .B(pi335), .C(pi079), .Y(po079));
  ADDER_G2_27_28_29 g159(.A(new_n928_), .B(pi335), .C(pi079), .Y(new_n930_));
  ADDER_G0_20_21    g160(.A(new_n930_), .B(pi336), .C(pi080), .Y(po080));
  ADDER_G2_27_28_29 g161(.A(new_n930_), .B(pi336), .C(pi080), .Y(new_n932_));
  ADDER_G0_20_21    g162(.A(new_n932_), .B(pi337), .C(pi081), .Y(po081));
  ADDER_G2_27_28_29 g163(.A(new_n932_), .B(pi337), .C(pi081), .Y(new_n934_));
  ADDER_G0_20_21    g164(.A(new_n934_), .B(pi338), .C(pi082), .Y(po082));
  ADDER_G2_27_28_29 g165(.A(new_n934_), .B(pi338), .C(pi082), .Y(new_n936_));
  ADDER_G0_20_21    g166(.A(new_n936_), .B(pi339), .C(pi083), .Y(po083));
  ADDER_G2_27_28_29 g167(.A(new_n936_), .B(pi339), .C(pi083), .Y(new_n938_));
  ADDER_G0_20_21    g168(.A(new_n938_), .B(pi340), .C(pi084), .Y(po084));
  ADDER_G2_27_28_29 g169(.A(new_n938_), .B(pi340), .C(pi084), .Y(new_n940_));
  ADDER_G0_20_21    g170(.A(new_n940_), .B(pi341), .C(pi085), .Y(po085));
  ADDER_G2_27_28_29 g171(.A(new_n940_), .B(pi341), .C(pi085), .Y(new_n942_));
  ADDER_G0_20_21    g172(.A(new_n942_), .B(pi342), .C(pi086), .Y(po086));
  ADDER_G2_27_28_29 g173(.A(new_n942_), .B(pi342), .C(pi086), .Y(new_n944_));
  ADDER_G0_20_21    g174(.A(new_n944_), .B(pi343), .C(pi087), .Y(po087));
  ADDER_G2_27_28_29 g175(.A(new_n944_), .B(pi343), .C(pi087), .Y(new_n946_));
  ADDER_G0_20_21    g176(.A(new_n946_), .B(pi344), .C(pi088), .Y(po088));
  ADDER_G2_27_28_29 g177(.A(new_n946_), .B(pi344), .C(pi088), .Y(new_n948_));
  ADDER_G0_20_21    g178(.A(new_n948_), .B(pi345), .C(pi089), .Y(po089));
  ADDER_G2_27_28_29 g179(.A(new_n948_), .B(pi345), .C(pi089), .Y(new_n950_));
  ADDER_G0_20_21    g180(.A(new_n950_), .B(pi346), .C(pi090), .Y(po090));
  ADDER_G2_27_28_29 g181(.A(new_n950_), .B(pi346), .C(pi090), .Y(new_n952_));
  ADDER_G0_20_21    g182(.A(new_n952_), .B(pi347), .C(pi091), .Y(po091));
  ADDER_G2_27_28_29 g183(.A(new_n952_), .B(pi347), .C(pi091), .Y(new_n954_));
  ADDER_G0_20_21    g184(.A(new_n954_), .B(pi348), .C(pi092), .Y(po092));
  ADDER_G2_27_28_29 g185(.A(new_n954_), .B(pi348), .C(pi092), .Y(new_n956_));
  ADDER_G0_20_21    g186(.A(new_n956_), .B(pi349), .C(pi093), .Y(po093));
  ADDER_G2_27_28_29 g187(.A(new_n956_), .B(pi349), .C(pi093), .Y(new_n958_));
  ADDER_G0_20_21    g188(.A(new_n958_), .B(pi350), .C(pi094), .Y(po094));
  ADDER_G2_27_28_29 g189(.A(new_n958_), .B(pi350), .C(pi094), .Y(new_n960_));
  ADDER_G0_20_21    g190(.A(new_n960_), .B(pi351), .C(pi095), .Y(po095));
  ADDER_G2_27_28_29 g191(.A(new_n960_), .B(pi351), .C(pi095), .Y(new_n962_));
  ADDER_G0_20_21    g192(.A(new_n962_), .B(pi352), .C(pi096), .Y(po096));
  ADDER_G2_27_28_29 g193(.A(new_n962_), .B(pi352), .C(pi096), .Y(new_n964_));
  ADDER_G0_20_21    g194(.A(new_n964_), .B(pi353), .C(pi097), .Y(po097));
  ADDER_G2_27_28_29 g195(.A(new_n964_), .B(pi353), .C(pi097), .Y(new_n966_));
  ADDER_G0_20_21    g196(.A(new_n966_), .B(pi354), .C(pi098), .Y(po098));
  ADDER_G2_27_28_29 g197(.A(new_n966_), .B(pi354), .C(pi098), .Y(new_n968_));
  ADDER_G0_20_21    g198(.A(new_n968_), .B(pi355), .C(pi099), .Y(po099));
  ADDER_G2_27_28_29 g199(.A(new_n968_), .B(pi355), .C(pi099), .Y(new_n970_));
  ADDER_G0_20_21    g200(.A(new_n970_), .B(pi356), .C(pi100), .Y(po100));
  ADDER_G2_27_28_29 g201(.A(new_n970_), .B(pi356), .C(pi100), .Y(new_n972_));
  ADDER_G0_20_21    g202(.A(new_n972_), .B(pi357), .C(pi101), .Y(po101));
  ADDER_G2_27_28_29 g203(.A(new_n972_), .B(pi357), .C(pi101), .Y(new_n974_));
  ADDER_G0_20_21    g204(.A(new_n974_), .B(pi358), .C(pi102), .Y(po102));
  ADDER_G2_27_28_29 g205(.A(new_n974_), .B(pi358), .C(pi102), .Y(new_n976_));
  ADDER_G0_20_21    g206(.A(new_n976_), .B(pi359), .C(pi103), .Y(po103));
  ADDER_G2_27_28_29 g207(.A(new_n976_), .B(pi359), .C(pi103), .Y(new_n978_));
  ADDER_G0_20_21    g208(.A(new_n978_), .B(pi360), .C(pi104), .Y(po104));
  ADDER_G2_27_28_29 g209(.A(new_n978_), .B(pi360), .C(pi104), .Y(new_n980_));
  ADDER_G0_20_21    g210(.A(new_n980_), .B(pi361), .C(pi105), .Y(po105));
  ADDER_G2_27_28_29 g211(.A(new_n980_), .B(pi361), .C(pi105), .Y(new_n982_));
  ADDER_G0_20_21    g212(.A(new_n982_), .B(pi362), .C(pi106), .Y(po106));
  ADDER_G2_27_28_29 g213(.A(new_n982_), .B(pi362), .C(pi106), .Y(new_n984_));
  ADDER_G0_20_21    g214(.A(new_n984_), .B(pi363), .C(pi107), .Y(po107));
  ADDER_G2_27_28_29 g215(.A(new_n984_), .B(pi363), .C(pi107), .Y(new_n986_));
  ADDER_G0_20_21    g216(.A(new_n986_), .B(pi364), .C(pi108), .Y(po108));
  ADDER_G2_27_28_29 g217(.A(new_n986_), .B(pi364), .C(pi108), .Y(new_n988_));
  ADDER_G0_20_21    g218(.A(new_n988_), .B(pi365), .C(pi109), .Y(po109));
  ADDER_G2_27_28_29 g219(.A(new_n988_), .B(pi365), .C(pi109), .Y(new_n990_));
  ADDER_G0_20_21    g220(.A(new_n990_), .B(pi366), .C(pi110), .Y(po110));
  ADDER_G2_27_28_29 g221(.A(new_n990_), .B(pi366), .C(pi110), .Y(new_n992_));
  ADDER_G0_20_21    g222(.A(new_n992_), .B(pi367), .C(pi111), .Y(po111));
  ADDER_G2_27_28_29 g223(.A(new_n992_), .B(pi367), .C(pi111), .Y(new_n994_));
  ADDER_G0_20_21    g224(.A(new_n994_), .B(pi368), .C(pi112), .Y(po112));
  ADDER_G2_27_28_29 g225(.A(new_n994_), .B(pi368), .C(pi112), .Y(new_n996_));
  ADDER_G0_20_21    g226(.A(new_n996_), .B(pi369), .C(pi113), .Y(po113));
  ADDER_G2_27_28_29 g227(.A(new_n996_), .B(pi369), .C(pi113), .Y(new_n998_));
  ADDER_G0_20_21    g228(.A(new_n998_), .B(pi370), .C(pi114), .Y(po114));
  ADDER_G2_27_28_29 g229(.A(new_n998_), .B(pi370), .C(pi114), .Y(new_n1000_));
  ADDER_G0_20_21    g230(.A(new_n1000_), .B(pi371), .C(pi115), .Y(po115));
  ADDER_G2_27_28_29 g231(.A(new_n1000_), .B(pi371), .C(pi115), .Y(new_n1002_));
  ADDER_G0_20_21    g232(.A(new_n1002_), .B(pi372), .C(pi116), .Y(po116));
  ADDER_G2_27_28_29 g233(.A(new_n1002_), .B(pi372), .C(pi116), .Y(new_n1004_));
  ADDER_G0_20_21    g234(.A(new_n1004_), .B(pi373), .C(pi117), .Y(po117));
  ADDER_G2_27_28_29 g235(.A(new_n1004_), .B(pi373), .C(pi117), .Y(new_n1006_));
  ADDER_G0_20_21    g236(.A(new_n1006_), .B(pi374), .C(pi118), .Y(po118));
  ADDER_G2_27_28_29 g237(.A(new_n1006_), .B(pi374), .C(pi118), .Y(new_n1008_));
  ADDER_G0_20_21    g238(.A(new_n1008_), .B(pi375), .C(pi119), .Y(po119));
  ADDER_G2_27_28_29 g239(.A(new_n1008_), .B(pi375), .C(pi119), .Y(new_n1010_));
  ADDER_G0_20_21    g240(.A(new_n1010_), .B(pi376), .C(pi120), .Y(po120));
  ADDER_G2_27_28_29 g241(.A(new_n1010_), .B(pi376), .C(pi120), .Y(new_n1012_));
  ADDER_G0_20_21    g242(.A(new_n1012_), .B(pi377), .C(pi121), .Y(po121));
  ADDER_G2_27_28_29 g243(.A(new_n1012_), .B(pi377), .C(pi121), .Y(new_n1014_));
  ADDER_G0_20_21    g244(.A(new_n1014_), .B(pi378), .C(pi122), .Y(po122));
  ADDER_G2_27_28_29 g245(.A(new_n1014_), .B(pi378), .C(pi122), .Y(new_n1016_));
  ADDER_G0_20_21    g246(.A(new_n1016_), .B(pi379), .C(pi123), .Y(po123));
  ADDER_G2_27_28_29 g247(.A(new_n1016_), .B(pi379), .C(pi123), .Y(new_n1018_));
  ADDER_G0_20_21    g248(.A(new_n1018_), .B(pi380), .C(pi124), .Y(po124));
  ADDER_G2_27_28_29 g249(.A(new_n1018_), .B(pi380), .C(pi124), .Y(new_n1020_));
  ADDER_G0_20_21    g250(.A(new_n1020_), .B(pi381), .C(pi125), .Y(po125));
  ADDER_G2_27_28_29 g251(.A(new_n1020_), .B(pi381), .C(pi125), .Y(new_n1022_));
  ADDER_G0_20_21    g252(.A(new_n1022_), .B(pi382), .C(pi126), .Y(po126));
  ADDER_G2_27_28_29 g253(.A(new_n1022_), .B(pi382), .C(pi126), .Y(new_n1024_));
  ADDER_G0_20_21    g254(.A(new_n1024_), .B(pi383), .C(pi127), .Y(po127));
  ADDER_G2_27_28_29 g255(.A(new_n1024_), .B(pi383), .C(pi127), .Y(new_n1026_));
  ADDER_G0_20_21    g256(.A(new_n1026_), .B(pi384), .C(pi128), .Y(po128));
  ADDER_G2_27_28_29 g257(.A(new_n1026_), .B(pi384), .C(pi128), .Y(new_n1028_));
  ADDER_G0_20_21    g258(.A(new_n1028_), .B(pi385), .C(pi129), .Y(po129));
  ADDER_G2_27_28_29 g259(.A(new_n1028_), .B(pi385), .C(pi129), .Y(new_n1030_));
  ADDER_G0_20_21    g260(.A(new_n1030_), .B(pi386), .C(pi130), .Y(po130));
  ADDER_G2_27_28_29 g261(.A(new_n1030_), .B(pi386), .C(pi130), .Y(new_n1032_));
  ADDER_G0_20_21    g262(.A(new_n1032_), .B(pi387), .C(pi131), .Y(po131));
  ADDER_G2_27_28_29 g263(.A(new_n1032_), .B(pi387), .C(pi131), .Y(new_n1034_));
  ADDER_G0_20_21    g264(.A(new_n1034_), .B(pi388), .C(pi132), .Y(po132));
  ADDER_G2_27_28_29 g265(.A(new_n1034_), .B(pi388), .C(pi132), .Y(new_n1036_));
  ADDER_G0_20_21    g266(.A(new_n1036_), .B(pi389), .C(pi133), .Y(po133));
  ADDER_G2_27_28_29 g267(.A(new_n1036_), .B(pi389), .C(pi133), .Y(new_n1038_));
  ADDER_G0_20_21    g268(.A(new_n1038_), .B(pi390), .C(pi134), .Y(po134));
  ADDER_G2_27_28_29 g269(.A(new_n1038_), .B(pi390), .C(pi134), .Y(new_n1040_));
  ADDER_G0_20_21    g270(.A(new_n1040_), .B(pi391), .C(pi135), .Y(po135));
  ADDER_G2_27_28_29 g271(.A(new_n1040_), .B(pi391), .C(pi135), .Y(new_n1042_));
  ADDER_G0_20_21    g272(.A(new_n1042_), .B(pi392), .C(pi136), .Y(po136));
  ADDER_G2_27_28_29 g273(.A(new_n1042_), .B(pi392), .C(pi136), .Y(new_n1044_));
  ADDER_G0_20_21    g274(.A(new_n1044_), .B(pi393), .C(pi137), .Y(po137));
  ADDER_G2_27_28_29 g275(.A(new_n1044_), .B(pi393), .C(pi137), .Y(new_n1046_));
  ADDER_G0_20_21    g276(.A(new_n1046_), .B(pi394), .C(pi138), .Y(po138));
  ADDER_G2_27_28_29 g277(.A(new_n1046_), .B(pi394), .C(pi138), .Y(new_n1048_));
  ADDER_G0_20_21    g278(.A(new_n1048_), .B(pi395), .C(pi139), .Y(po139));
  ADDER_G2_27_28_29 g279(.A(new_n1048_), .B(pi395), .C(pi139), .Y(new_n1050_));
  ADDER_G0_20_21    g280(.A(new_n1050_), .B(pi396), .C(pi140), .Y(po140));
  ADDER_G2_27_28_29 g281(.A(new_n1050_), .B(pi396), .C(pi140), .Y(new_n1052_));
  ADDER_G0_20_21    g282(.A(new_n1052_), .B(pi397), .C(pi141), .Y(po141));
  ADDER_G2_27_28_29 g283(.A(new_n1052_), .B(pi397), .C(pi141), .Y(new_n1054_));
  ADDER_G0_20_21    g284(.A(new_n1054_), .B(pi398), .C(pi142), .Y(po142));
  ADDER_G2_27_28_29 g285(.A(new_n1054_), .B(pi398), .C(pi142), .Y(new_n1056_));
  ADDER_G0_20_21    g286(.A(new_n1056_), .B(pi399), .C(pi143), .Y(po143));
  ADDER_G2_27_28_29 g287(.A(new_n1056_), .B(pi399), .C(pi143), .Y(new_n1058_));
  ADDER_G0_20_21    g288(.A(new_n1058_), .B(pi400), .C(pi144), .Y(po144));
  ADDER_G2_27_28_29 g289(.A(new_n1058_), .B(pi400), .C(pi144), .Y(new_n1060_));
  ADDER_G0_20_21    g290(.A(new_n1060_), .B(pi401), .C(pi145), .Y(po145));
  ADDER_G2_27_28_29 g291(.A(new_n1060_), .B(pi401), .C(pi145), .Y(new_n1062_));
  ADDER_G0_20_21    g292(.A(new_n1062_), .B(pi402), .C(pi146), .Y(po146));
  ADDER_G2_27_28_29 g293(.A(new_n1062_), .B(pi402), .C(pi146), .Y(new_n1064_));
  ADDER_G0_20_21    g294(.A(new_n1064_), .B(pi403), .C(pi147), .Y(po147));
  ADDER_G2_27_28_29 g295(.A(new_n1064_), .B(pi403), .C(pi147), .Y(new_n1066_));
  ADDER_G0_20_21    g296(.A(new_n1066_), .B(pi404), .C(pi148), .Y(po148));
  ADDER_G2_27_28_29 g297(.A(new_n1066_), .B(pi404), .C(pi148), .Y(new_n1068_));
  ADDER_G0_20_21    g298(.A(new_n1068_), .B(pi405), .C(pi149), .Y(po149));
  ADDER_G2_27_28_29 g299(.A(new_n1068_), .B(pi405), .C(pi149), .Y(new_n1070_));
  ADDER_G0_20_21    g300(.A(new_n1070_), .B(pi406), .C(pi150), .Y(po150));
  ADDER_G2_27_28_29 g301(.A(new_n1070_), .B(pi406), .C(pi150), .Y(new_n1072_));
  ADDER_G0_20_21    g302(.A(new_n1072_), .B(pi407), .C(pi151), .Y(po151));
  ADDER_G2_27_28_29 g303(.A(new_n1072_), .B(pi407), .C(pi151), .Y(new_n1074_));
  ADDER_G0_20_21    g304(.A(new_n1074_), .B(pi408), .C(pi152), .Y(po152));
  ADDER_G2_27_28_29 g305(.A(new_n1074_), .B(pi408), .C(pi152), .Y(new_n1076_));
  ADDER_G0_20_21    g306(.A(new_n1076_), .B(pi409), .C(pi153), .Y(po153));
  ADDER_G2_27_28_29 g307(.A(new_n1076_), .B(pi409), .C(pi153), .Y(new_n1078_));
  ADDER_G0_20_21    g308(.A(new_n1078_), .B(pi410), .C(pi154), .Y(po154));
  ADDER_G2_27_28_29 g309(.A(new_n1078_), .B(pi410), .C(pi154), .Y(new_n1080_));
  ADDER_G0_20_21    g310(.A(new_n1080_), .B(pi411), .C(pi155), .Y(po155));
  ADDER_G2_27_28_29 g311(.A(new_n1080_), .B(pi411), .C(pi155), .Y(new_n1082_));
  ADDER_G0_20_21    g312(.A(new_n1082_), .B(pi412), .C(pi156), .Y(po156));
  ADDER_G2_27_28_29 g313(.A(new_n1082_), .B(pi412), .C(pi156), .Y(new_n1084_));
  ADDER_G0_20_21    g314(.A(new_n1084_), .B(pi413), .C(pi157), .Y(po157));
  ADDER_G2_27_28_29 g315(.A(new_n1084_), .B(pi413), .C(pi157), .Y(new_n1086_));
  ADDER_G0_20_21    g316(.A(new_n1086_), .B(pi414), .C(pi158), .Y(po158));
  ADDER_G2_27_28_29 g317(.A(new_n1086_), .B(pi414), .C(pi158), .Y(new_n1088_));
  ADDER_G0_20_21    g318(.A(new_n1088_), .B(pi415), .C(pi159), .Y(po159));
  ADDER_G2_27_28_29 g319(.A(new_n1088_), .B(pi415), .C(pi159), .Y(new_n1090_));
  ADDER_G0_20_21    g320(.A(new_n1090_), .B(pi416), .C(pi160), .Y(po160));
  ADDER_G2_27_28_29 g321(.A(new_n1090_), .B(pi416), .C(pi160), .Y(new_n1092_));
  ADDER_G0_20_21    g322(.A(new_n1092_), .B(pi417), .C(pi161), .Y(po161));
  ADDER_G2_27_28_29 g323(.A(new_n1092_), .B(pi417), .C(pi161), .Y(new_n1094_));
  ADDER_G0_20_21    g324(.A(new_n1094_), .B(pi418), .C(pi162), .Y(po162));
  ADDER_G2_27_28_29 g325(.A(new_n1094_), .B(pi418), .C(pi162), .Y(new_n1096_));
  ADDER_G0_20_21    g326(.A(new_n1096_), .B(pi419), .C(pi163), .Y(po163));
  ADDER_G2_27_28_29 g327(.A(new_n1096_), .B(pi419), .C(pi163), .Y(new_n1098_));
  ADDER_G0_20_21    g328(.A(new_n1098_), .B(pi420), .C(pi164), .Y(po164));
  ADDER_G2_27_28_29 g329(.A(new_n1098_), .B(pi420), .C(pi164), .Y(new_n1100_));
  ADDER_G0_20_21    g330(.A(new_n1100_), .B(pi421), .C(pi165), .Y(po165));
  ADDER_G2_27_28_29 g331(.A(new_n1100_), .B(pi421), .C(pi165), .Y(new_n1102_));
  ADDER_G0_20_21    g332(.A(new_n1102_), .B(pi422), .C(pi166), .Y(po166));
  ADDER_G2_27_28_29 g333(.A(new_n1102_), .B(pi422), .C(pi166), .Y(new_n1104_));
  ADDER_G0_20_21    g334(.A(new_n1104_), .B(pi423), .C(pi167), .Y(po167));
  ADDER_G2_27_28_29 g335(.A(new_n1104_), .B(pi423), .C(pi167), .Y(new_n1106_));
  ADDER_G0_20_21    g336(.A(new_n1106_), .B(pi424), .C(pi168), .Y(po168));
  ADDER_G2_27_28_29 g337(.A(new_n1106_), .B(pi424), .C(pi168), .Y(new_n1108_));
  ADDER_G0_20_21    g338(.A(new_n1108_), .B(pi425), .C(pi169), .Y(po169));
  ADDER_G2_27_28_29 g339(.A(new_n1108_), .B(pi425), .C(pi169), .Y(new_n1110_));
  ADDER_G0_20_21    g340(.A(new_n1110_), .B(pi426), .C(pi170), .Y(po170));
  ADDER_G2_27_28_29 g341(.A(new_n1110_), .B(pi426), .C(pi170), .Y(new_n1112_));
  ADDER_G0_20_21    g342(.A(new_n1112_), .B(pi427), .C(pi171), .Y(po171));
  ADDER_G2_27_28_29 g343(.A(new_n1112_), .B(pi427), .C(pi171), .Y(new_n1114_));
  ADDER_G0_20_21    g344(.A(new_n1114_), .B(pi428), .C(pi172), .Y(po172));
  ADDER_G2_27_28_29 g345(.A(new_n1114_), .B(pi428), .C(pi172), .Y(new_n1116_));
  ADDER_G0_20_21    g346(.A(new_n1116_), .B(pi429), .C(pi173), .Y(po173));
  ADDER_G2_27_28_29 g347(.A(new_n1116_), .B(pi429), .C(pi173), .Y(new_n1118_));
  ADDER_G0_20_21    g348(.A(new_n1118_), .B(pi430), .C(pi174), .Y(po174));
  ADDER_G2_27_28_29 g349(.A(new_n1118_), .B(pi430), .C(pi174), .Y(new_n1120_));
  ADDER_G0_20_21    g350(.A(new_n1120_), .B(pi431), .C(pi175), .Y(po175));
  ADDER_G2_27_28_29 g351(.A(new_n1120_), .B(pi431), .C(pi175), .Y(new_n1122_));
  ADDER_G0_20_21    g352(.A(new_n1122_), .B(pi432), .C(pi176), .Y(po176));
  ADDER_G2_27_28_29 g353(.A(new_n1122_), .B(pi432), .C(pi176), .Y(new_n1124_));
  ADDER_G0_20_21    g354(.A(new_n1124_), .B(pi433), .C(pi177), .Y(po177));
  ADDER_G2_27_28_29 g355(.A(new_n1124_), .B(pi433), .C(pi177), .Y(new_n1126_));
  ADDER_G0_20_21    g356(.A(new_n1126_), .B(pi434), .C(pi178), .Y(po178));
  ADDER_G2_27_28_29 g357(.A(new_n1126_), .B(pi434), .C(pi178), .Y(new_n1128_));
  ADDER_G0_20_21    g358(.A(new_n1128_), .B(pi435), .C(pi179), .Y(po179));
  ADDER_G2_27_28_29 g359(.A(new_n1128_), .B(pi435), .C(pi179), .Y(new_n1130_));
  ADDER_G0_20_21    g360(.A(new_n1130_), .B(pi436), .C(pi180), .Y(po180));
  ADDER_G2_27_28_29 g361(.A(new_n1130_), .B(pi436), .C(pi180), .Y(new_n1132_));
  ADDER_G0_20_21    g362(.A(new_n1132_), .B(pi437), .C(pi181), .Y(po181));
  ADDER_G2_27_28_29 g363(.A(new_n1132_), .B(pi437), .C(pi181), .Y(new_n1134_));
  ADDER_G0_20_21    g364(.A(new_n1134_), .B(pi438), .C(pi182), .Y(po182));
  ADDER_G2_27_28_29 g365(.A(new_n1134_), .B(pi438), .C(pi182), .Y(new_n1136_));
  ADDER_G0_20_21    g366(.A(new_n1136_), .B(pi439), .C(pi183), .Y(po183));
  ADDER_G2_27_28_29 g367(.A(new_n1136_), .B(pi439), .C(pi183), .Y(new_n1138_));
  ADDER_G0_20_21    g368(.A(new_n1138_), .B(pi440), .C(pi184), .Y(po184));
  ADDER_G2_27_28_29 g369(.A(new_n1138_), .B(pi440), .C(pi184), .Y(new_n1140_));
  ADDER_G0_20_21    g370(.A(new_n1140_), .B(pi441), .C(pi185), .Y(po185));
  ADDER_G2_27_28_29 g371(.A(new_n1140_), .B(pi441), .C(pi185), .Y(new_n1142_));
  ADDER_G0_20_21    g372(.A(new_n1142_), .B(pi442), .C(pi186), .Y(po186));
  ADDER_G2_27_28_29 g373(.A(new_n1142_), .B(pi442), .C(pi186), .Y(new_n1144_));
  ADDER_G0_20_21    g374(.A(new_n1144_), .B(pi443), .C(pi187), .Y(po187));
  ADDER_G2_27_28_29 g375(.A(new_n1144_), .B(pi443), .C(pi187), .Y(new_n1146_));
  ADDER_G0_20_21    g376(.A(new_n1146_), .B(pi444), .C(pi188), .Y(po188));
  ADDER_G2_27_28_29 g377(.A(new_n1146_), .B(pi444), .C(pi188), .Y(new_n1148_));
  ADDER_G0_20_21    g378(.A(new_n1148_), .B(pi445), .C(pi189), .Y(po189));
  ADDER_G2_27_28_29 g379(.A(new_n1148_), .B(pi445), .C(pi189), .Y(new_n1150_));
  ADDER_G0_20_21    g380(.A(new_n1150_), .B(pi446), .C(pi190), .Y(po190));
  ADDER_G2_27_28_29 g381(.A(new_n1150_), .B(pi446), .C(pi190), .Y(new_n1152_));
  ADDER_G0_20_21    g382(.A(new_n1152_), .B(pi447), .C(pi191), .Y(po191));
  ADDER_G2_27_28_29 g383(.A(new_n1152_), .B(pi447), .C(pi191), .Y(new_n1154_));
  ADDER_G0_20_21    g384(.A(new_n1154_), .B(pi448), .C(pi192), .Y(po192));
  ADDER_G2_27_28_29 g385(.A(new_n1154_), .B(pi448), .C(pi192), .Y(new_n1156_));
  ADDER_G0_20_21    g386(.A(new_n1156_), .B(pi449), .C(pi193), .Y(po193));
  ADDER_G2_27_28_29 g387(.A(new_n1156_), .B(pi449), .C(pi193), .Y(new_n1158_));
  ADDER_G0_20_21    g388(.A(new_n1158_), .B(pi450), .C(pi194), .Y(po194));
  ADDER_G2_27_28_29 g389(.A(new_n1158_), .B(pi450), .C(pi194), .Y(new_n1160_));
  ADDER_G0_20_21    g390(.A(new_n1160_), .B(pi451), .C(pi195), .Y(po195));
  ADDER_G2_27_28_29 g391(.A(new_n1160_), .B(pi451), .C(pi195), .Y(new_n1162_));
  ADDER_G0_20_21    g392(.A(new_n1162_), .B(pi452), .C(pi196), .Y(po196));
  ADDER_G2_27_28_29 g393(.A(new_n1162_), .B(pi452), .C(pi196), .Y(new_n1164_));
  ADDER_G0_20_21    g394(.A(new_n1164_), .B(pi453), .C(pi197), .Y(po197));
  ADDER_G2_27_28_29 g395(.A(new_n1164_), .B(pi453), .C(pi197), .Y(new_n1166_));
  ADDER_G0_20_21    g396(.A(new_n1166_), .B(pi454), .C(pi198), .Y(po198));
  ADDER_G2_27_28_29 g397(.A(new_n1166_), .B(pi454), .C(pi198), .Y(new_n1168_));
  ADDER_G0_20_21    g398(.A(new_n1168_), .B(pi455), .C(pi199), .Y(po199));
  ADDER_G2_27_28_29 g399(.A(new_n1168_), .B(pi455), .C(pi199), .Y(new_n1170_));
  ADDER_G0_20_21    g400(.A(new_n1170_), .B(pi456), .C(pi200), .Y(po200));
  ADDER_G2_27_28_29 g401(.A(new_n1170_), .B(pi456), .C(pi200), .Y(new_n1172_));
  ADDER_G0_20_21    g402(.A(new_n1172_), .B(pi457), .C(pi201), .Y(po201));
  ADDER_G2_27_28_29 g403(.A(new_n1172_), .B(pi457), .C(pi201), .Y(new_n1174_));
  ADDER_G0_20_21    g404(.A(new_n1174_), .B(pi458), .C(pi202), .Y(po202));
  ADDER_G2_27_28_29 g405(.A(new_n1174_), .B(pi458), .C(pi202), .Y(new_n1176_));
  ADDER_G0_20_21    g406(.A(new_n1176_), .B(pi459), .C(pi203), .Y(po203));
  ADDER_G2_27_28_29 g407(.A(new_n1176_), .B(pi459), .C(pi203), .Y(new_n1178_));
  ADDER_G0_20_21    g408(.A(new_n1178_), .B(pi460), .C(pi204), .Y(po204));
  ADDER_G2_27_28_29 g409(.A(new_n1178_), .B(pi460), .C(pi204), .Y(new_n1180_));
  ADDER_G0_20_21    g410(.A(new_n1180_), .B(pi461), .C(pi205), .Y(po205));
  ADDER_G2_27_28_29 g411(.A(new_n1180_), .B(pi461), .C(pi205), .Y(new_n1182_));
  ADDER_G0_20_21    g412(.A(new_n1182_), .B(pi462), .C(pi206), .Y(po206));
  ADDER_G2_27_28_29 g413(.A(new_n1182_), .B(pi462), .C(pi206), .Y(new_n1184_));
  ADDER_G0_20_21    g414(.A(new_n1184_), .B(pi463), .C(pi207), .Y(po207));
  ADDER_G2_27_28_29 g415(.A(new_n1184_), .B(pi463), .C(pi207), .Y(new_n1186_));
  ADDER_G0_20_21    g416(.A(new_n1186_), .B(pi464), .C(pi208), .Y(po208));
  ADDER_G2_27_28_29 g417(.A(new_n1186_), .B(pi464), .C(pi208), .Y(new_n1188_));
  ADDER_G0_20_21    g418(.A(new_n1188_), .B(pi465), .C(pi209), .Y(po209));
  ADDER_G2_27_28_29 g419(.A(new_n1188_), .B(pi465), .C(pi209), .Y(new_n1190_));
  ADDER_G0_20_21    g420(.A(new_n1190_), .B(pi466), .C(pi210), .Y(po210));
  ADDER_G2_27_28_29 g421(.A(new_n1190_), .B(pi466), .C(pi210), .Y(new_n1192_));
  ADDER_G0_20_21    g422(.A(new_n1192_), .B(pi467), .C(pi211), .Y(po211));
  ADDER_G2_27_28_29 g423(.A(new_n1192_), .B(pi467), .C(pi211), .Y(new_n1194_));
  ADDER_G0_20_21    g424(.A(new_n1194_), .B(pi468), .C(pi212), .Y(po212));
  ADDER_G2_27_28_29 g425(.A(new_n1194_), .B(pi468), .C(pi212), .Y(new_n1196_));
  ADDER_G0_20_21    g426(.A(new_n1196_), .B(pi469), .C(pi213), .Y(po213));
  ADDER_G2_27_28_29 g427(.A(new_n1196_), .B(pi469), .C(pi213), .Y(new_n1198_));
  ADDER_G0_20_21    g428(.A(new_n1198_), .B(pi470), .C(pi214), .Y(po214));
  ADDER_G2_27_28_29 g429(.A(new_n1198_), .B(pi470), .C(pi214), .Y(new_n1200_));
  ADDER_G0_20_21    g430(.A(new_n1200_), .B(pi471), .C(pi215), .Y(po215));
  ADDER_G2_27_28_29 g431(.A(new_n1200_), .B(pi471), .C(pi215), .Y(new_n1202_));
  ADDER_G0_20_21    g432(.A(new_n1202_), .B(pi472), .C(pi216), .Y(po216));
  ADDER_G2_27_28_29 g433(.A(new_n1202_), .B(pi472), .C(pi216), .Y(new_n1204_));
  ADDER_G0_20_21    g434(.A(new_n1204_), .B(pi473), .C(pi217), .Y(po217));
  ADDER_G2_27_28_29 g435(.A(new_n1204_), .B(pi473), .C(pi217), .Y(new_n1206_));
  ADDER_G0_20_21    g436(.A(new_n1206_), .B(pi474), .C(pi218), .Y(po218));
  ADDER_G2_27_28_29 g437(.A(new_n1206_), .B(pi474), .C(pi218), .Y(new_n1208_));
  ADDER_G0_20_21    g438(.A(new_n1208_), .B(pi475), .C(pi219), .Y(po219));
  ADDER_G2_27_28_29 g439(.A(new_n1208_), .B(pi475), .C(pi219), .Y(new_n1210_));
  ADDER_G0_20_21    g440(.A(new_n1210_), .B(pi476), .C(pi220), .Y(po220));
  ADDER_G2_27_28_29 g441(.A(new_n1210_), .B(pi476), .C(pi220), .Y(new_n1212_));
  ADDER_G0_20_21    g442(.A(new_n1212_), .B(pi477), .C(pi221), .Y(po221));
  ADDER_G2_27_28_29 g443(.A(new_n1212_), .B(pi477), .C(pi221), .Y(new_n1214_));
  ADDER_G0_20_21    g444(.A(new_n1214_), .B(pi478), .C(pi222), .Y(po222));
  ADDER_G2_27_28_29 g445(.A(new_n1214_), .B(pi478), .C(pi222), .Y(new_n1216_));
  ADDER_G0_20_21    g446(.A(new_n1216_), .B(pi479), .C(pi223), .Y(po223));
  ADDER_G2_27_28_29 g447(.A(new_n1216_), .B(pi479), .C(pi223), .Y(new_n1218_));
  ADDER_G0_20_21    g448(.A(new_n1218_), .B(pi480), .C(pi224), .Y(po224));
  ADDER_G2_27_28_29 g449(.A(new_n1218_), .B(pi480), .C(pi224), .Y(new_n1220_));
  ADDER_G0_20_21    g450(.A(new_n1220_), .B(pi481), .C(pi225), .Y(po225));
  ADDER_G2_27_28_29 g451(.A(new_n1220_), .B(pi481), .C(pi225), .Y(new_n1222_));
  ADDER_G0_20_21    g452(.A(new_n1222_), .B(pi482), .C(pi226), .Y(po226));
  ADDER_G2_27_28_29 g453(.A(new_n1222_), .B(pi482), .C(pi226), .Y(new_n1224_));
  ADDER_G0_20_21    g454(.A(new_n1224_), .B(pi483), .C(pi227), .Y(po227));
  ADDER_G2_27_28_29 g455(.A(new_n1224_), .B(pi483), .C(pi227), .Y(new_n1226_));
  ADDER_G0_20_21    g456(.A(new_n1226_), .B(pi484), .C(pi228), .Y(po228));
  ADDER_G2_27_28_29 g457(.A(new_n1226_), .B(pi484), .C(pi228), .Y(new_n1228_));
  ADDER_G0_20_21    g458(.A(new_n1228_), .B(pi485), .C(pi229), .Y(po229));
  ADDER_G2_27_28_29 g459(.A(new_n1228_), .B(pi485), .C(pi229), .Y(new_n1230_));
  ADDER_G0_20_21    g460(.A(new_n1230_), .B(pi486), .C(pi230), .Y(po230));
  ADDER_G2_27_28_29 g461(.A(new_n1230_), .B(pi486), .C(pi230), .Y(new_n1232_));
  ADDER_G0_20_21    g462(.A(new_n1232_), .B(pi487), .C(pi231), .Y(po231));
  ADDER_G2_27_28_29 g463(.A(new_n1232_), .B(pi487), .C(pi231), .Y(new_n1234_));
  ADDER_G0_20_21    g464(.A(new_n1234_), .B(pi488), .C(pi232), .Y(po232));
  ADDER_G2_27_28_29 g465(.A(new_n1234_), .B(pi488), .C(pi232), .Y(new_n1236_));
  ADDER_G0_20_21    g466(.A(new_n1236_), .B(pi489), .C(pi233), .Y(po233));
  ADDER_G2_27_28_29 g467(.A(new_n1236_), .B(pi489), .C(pi233), .Y(new_n1238_));
  ADDER_G0_20_21    g468(.A(new_n1238_), .B(pi490), .C(pi234), .Y(po234));
  ADDER_G2_27_28_29 g469(.A(new_n1238_), .B(pi490), .C(pi234), .Y(new_n1240_));
  ADDER_G0_20_21    g470(.A(new_n1240_), .B(pi491), .C(pi235), .Y(po235));
  ADDER_G2_27_28_29 g471(.A(new_n1240_), .B(pi491), .C(pi235), .Y(new_n1242_));
  ADDER_G0_20_21    g472(.A(new_n1242_), .B(pi492), .C(pi236), .Y(po236));
  ADDER_G2_27_28_29 g473(.A(new_n1242_), .B(pi492), .C(pi236), .Y(new_n1244_));
  ADDER_G0_20_21    g474(.A(new_n1244_), .B(pi493), .C(pi237), .Y(po237));
  ADDER_G2_27_28_29 g475(.A(new_n1244_), .B(pi493), .C(pi237), .Y(new_n1246_));
  ADDER_G0_20_21    g476(.A(new_n1246_), .B(pi494), .C(pi238), .Y(po238));
  ADDER_G2_27_28_29 g477(.A(new_n1246_), .B(pi494), .C(pi238), .Y(new_n1248_));
  ADDER_G0_20_21    g478(.A(new_n1248_), .B(pi495), .C(pi239), .Y(po239));
  ADDER_G2_27_28_29 g479(.A(new_n1248_), .B(pi495), .C(pi239), .Y(new_n1250_));
  ADDER_G0_20_21    g480(.A(new_n1250_), .B(pi496), .C(pi240), .Y(po240));
  ADDER_G2_27_28_29 g481(.A(new_n1250_), .B(pi496), .C(pi240), .Y(new_n1252_));
  ADDER_G0_20_21    g482(.A(new_n1252_), .B(pi497), .C(pi241), .Y(po241));
  ADDER_G2_27_28_29 g483(.A(new_n1252_), .B(pi497), .C(pi241), .Y(new_n1254_));
  ADDER_G0_20_21    g484(.A(new_n1254_), .B(pi498), .C(pi242), .Y(po242));
  ADDER_G2_27_28_29 g485(.A(new_n1254_), .B(pi498), .C(pi242), .Y(new_n1256_));
  ADDER_G0_20_21    g486(.A(new_n1256_), .B(pi499), .C(pi243), .Y(po243));
  ADDER_G2_27_28_29 g487(.A(new_n1256_), .B(pi499), .C(pi243), .Y(new_n1258_));
  ADDER_G0_20_21    g488(.A(new_n1258_), .B(pi500), .C(pi244), .Y(po244));
  ADDER_G2_27_28_29 g489(.A(new_n1258_), .B(pi500), .C(pi244), .Y(new_n1260_));
  ADDER_G0_20_21    g490(.A(new_n1260_), .B(pi501), .C(pi245), .Y(po245));
  ADDER_G2_27_28_29 g491(.A(new_n1260_), .B(pi501), .C(pi245), .Y(new_n1262_));
  ADDER_G0_20_21    g492(.A(new_n1262_), .B(pi502), .C(pi246), .Y(po246));
  ADDER_G2_27_28_29 g493(.A(new_n1262_), .B(pi502), .C(pi246), .Y(new_n1264_));
  ADDER_G0_20_21    g494(.A(new_n1264_), .B(pi503), .C(pi247), .Y(po247));
  ADDER_G2_27_28_29 g495(.A(new_n1264_), .B(pi503), .C(pi247), .Y(new_n1266_));
  ADDER_G0_20_21    g496(.A(new_n1266_), .B(pi504), .C(pi248), .Y(po248));
  ADDER_G2_27_28_29 g497(.A(new_n1266_), .B(pi504), .C(pi248), .Y(new_n1268_));
  ADDER_G0_20_21    g498(.A(new_n1268_), .B(pi505), .C(pi249), .Y(po249));
  ADDER_G2_27_28_29 g499(.A(new_n1268_), .B(pi505), .C(pi249), .Y(new_n1270_));
  ADDER_G0_20_21    g500(.A(new_n1270_), .B(pi506), .C(pi250), .Y(po250));
  ADDER_G2_27_28_29 g501(.A(new_n1270_), .B(pi506), .C(pi250), .Y(new_n1272_));
  ADDER_G0_20_21    g502(.A(new_n1272_), .B(pi507), .C(pi251), .Y(po251));
  ADDER_G2_27_28_29 g503(.A(new_n1272_), .B(pi507), .C(pi251), .Y(new_n1274_));
  ADDER_G0_20_21    g504(.A(new_n1274_), .B(pi508), .C(pi252), .Y(po252));
  ADDER_G2_27_28_29 g505(.A(new_n1274_), .B(pi508), .C(pi252), .Y(new_n1276_));
  ADDER_G0_20_21    g506(.A(new_n1276_), .B(pi509), .C(pi253), .Y(po253));
  ADDER_G2_27_28_29 g507(.A(new_n1276_), .B(pi509), .C(pi253), .Y(new_n1278_));
  ADDER_G0_20_21    g508(.A(new_n1278_), .B(pi510), .C(pi254), .Y(po254));
  ADDER_G2_27_28_29 g509(.A(new_n1278_), .B(pi510), .C(pi254), .Y(new_n1280_));
  ADDER_G0_20_21    g510(.A(new_n1280_), .B(pi511), .C(pi255), .Y(po255));
  ADDER_G2_27_28_29 g511(.A(new_n1280_), .B(pi511), .C(pi255), .Y(po256));
endmodule


