.SUBCKT ROUTER_G1_38_39 A B C Y VCC GND
MclCO34LK_0#0 clCO34LK_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_0#1 VCC B clCO34LK_0#Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_0#2 clCO34LK_0#a_9_6# C GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_0#3 clCO34LK_0#Y B clCO34LK_0#a_9_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_1#0 Y clCO34LK_0#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_1#1 VCC A Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_1#2 clCO34LK_1#a_9_6# clCO34LK_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCO34LK_1#3 Y A clCO34LK_1#a_9_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 2|3|NAND2X1|NAND2X1=1|INPUT:Y-NAND2X1:A,B=3|NAND2X1:Y-NAND2X1:A,B=1|11101
* 18 occurrences in design
* each contains 2 cells
* pin map: {'x13': 'A', 'n106': 'B', 'n68': 'C'} {'n147': 'Y'}
* function: ~A|(B&C)
* Example occurence:
*   .subckt NAND2X1 A=n68 B=n106 Y=n107
*   .subckt NAND2X1 A=n107 B=x13 Y=n147
