.SUBCKT BAR_G3_0_2 A B C VDD VSS Y
MclWT24XJ_0#M0 clWT24XJ_0#Y C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_0#M1 clWT24XJ_0#Y C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_1#cl0S5SEU_0#M3 clWT24XJ_1#cl0S5SEU_0#net16 A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MclWT24XJ_1#cl0S5SEU_0#M2 clWT24XJ_1#cl0S5SEU_0#Y clWT24XJ_0#Y clWT24XJ_1#cl0S5SEU_0#net16 VSS nmos_lvt w=162.00n l=20n nfin=6
MclWT24XJ_1#cl0S5SEU_0#M1 clWT24XJ_1#cl0S5SEU_0#Y clWT24XJ_0#Y VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_1#cl0S5SEU_0#M0 clWT24XJ_1#cl0S5SEU_0#Y A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#M5 VSS clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net7 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#Y VSS nmos_lvt w=162.00n l=20n nfin=6
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#M1 VSS clWT24XJ_1#cl0S5SEU_1#C clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#M2 VSS B clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#M0 VDD clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net7 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#Y VDD pmos_lvt w=162.00n l=20n nfin=6
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#M4 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net15 clWT24XJ_1#cl0S5SEU_1#C clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net7 VDD pmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#M3 VDD B clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#net15 VDD pmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#M4 Y clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net10 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#M1 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net10 clWT24XJ_1#cl0S5SEU_0#Y VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#M0 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net10 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#Y VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#M5 Y clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net10 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#M3 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net20 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_0#Y VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MclWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#M2 clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net10 clWT24XJ_1#cl0S5SEU_0#Y clWT24XJ_1#cl0S5SEU_1#clB6EYAY_1#net20 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS 
* pattern code: 4|3|BAR_G2_3_5|INVx1=1|INPUT:Y-BAR_G2_3_5:A=1|INPUT:Y-BAR_G2_3_5:C=1|INPUT:Y-INVx1:A=1|INVx1:Y-BAR_G2_3_5:B=1|01111
* 408 occurrences in design
* each contains 2 cells
* function: (B&C)|(~A&~C)
* Example occurence:
*   .subckt INVx1 A=x128 Y=n250
*   .subckt BAR_G2_3_5 A=x57 B=n250 C=n188 Y=n358
