.SUBCKT SQRT_G0_173_198_231_260 A B C Y VCC GND
MclA3G2L7_0#0 VCC B clA3G2L7_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#1 clA3G2L7_0#a_18_54# clA3G2L7_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#2 clA3G2L7_0#Y clA3G2L7_0#a_2_6# clA3G2L7_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#3 clA3G2L7_0#a_35_54# B clA3G2L7_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#4 VCC C clA3G2L7_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#5 clA3G2L7_0#a_12_41# C VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#6 GND B clA3G2L7_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#7 clA3G2L7_0#a_18_6# clA3G2L7_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#8 clA3G2L7_0#Y B clA3G2L7_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#9 clA3G2L7_0#a_35_6# clA3G2L7_0#a_2_6# clA3G2L7_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#10 GND C clA3G2L7_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_0#11 clA3G2L7_0#a_12_41# C GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_1#0 clA3G2L7_1#Y clA3G2L7_0#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_1#1 clA3G2L7_1#Y clA3G2L7_0#Y GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#0 VCC A clA3G2L7_2#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#1 clA3G2L7_2#a_18_54# clA3G2L7_2#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#2 clA3G2L7_2#Y clA3G2L7_2#a_2_6# clA3G2L7_2#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#3 clA3G2L7_2#a_35_54# A clA3G2L7_2#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#4 VCC clA3G2L7_1#Y clA3G2L7_2#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#5 clA3G2L7_2#a_12_41# clA3G2L7_1#Y VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#6 GND A clA3G2L7_2#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#7 clA3G2L7_2#a_18_6# clA3G2L7_2#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#8 clA3G2L7_2#Y A clA3G2L7_2#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#9 clA3G2L7_2#a_35_6# clA3G2L7_2#a_2_6# clA3G2L7_2#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#10 GND clA3G2L7_1#Y clA3G2L7_2#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_2#11 clA3G2L7_2#a_12_41# clA3G2L7_1#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_3#0 Y clA3G2L7_2#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclA3G2L7_3#1 Y clA3G2L7_2#Y GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 4|3|INVX1|INVX1=1|XNOR2X1=2|INPUT:Y-XNOR2X1:A,B=3|INVX1:Y-XNOR2X1:A,B=1|XNOR2X1:Y-INVX1:A=2|1110111
* 1451 occurrences in design
* each contains 4 cells
* pin map: {'n488': 'A', 'n417': 'B', 'n350': 'C'} {'n490': 'Y'}
* function: (A&B&C)|(A&~B&~C)|(B&~A&~C)|(C&~A&~B)
* Example occurence:
*   .subckt XNOR2X1 A=n417 B=n350 Y=n418
*   .subckt INVX1 A=n418 Y=n419
*   .subckt XNOR2X1 A=n488 B=n419 Y=n489
*   .subckt INVX1 A=n489 Y=n490
