.SUBCKT VOTER_G3_6_8 A B C D Y VCC GND
MclAEAKO2_0#clCZWK1K_0#0 VCC C clAEAKO2_0#clCZWK1K_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#1 clAEAKO2_0#clCZWK1K_0#a_18_54# clAEAKO2_0#clCZWK1K_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#2 clAEAKO2_0#clCZWK1K_0#Y clAEAKO2_0#clCZWK1K_0#a_2_6# clAEAKO2_0#clCZWK1K_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#3 clAEAKO2_0#clCZWK1K_0#a_35_54# C clAEAKO2_0#clCZWK1K_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#4 VCC D clAEAKO2_0#clCZWK1K_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#5 clAEAKO2_0#clCZWK1K_0#a_12_41# D VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#6 GND C clAEAKO2_0#clCZWK1K_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#7 clAEAKO2_0#clCZWK1K_0#a_18_6# clAEAKO2_0#clCZWK1K_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#8 clAEAKO2_0#clCZWK1K_0#Y C clAEAKO2_0#clCZWK1K_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#9 clAEAKO2_0#clCZWK1K_0#a_35_6# clAEAKO2_0#clCZWK1K_0#a_2_6# clAEAKO2_0#clCZWK1K_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#10 GND D clAEAKO2_0#clCZWK1K_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_0#11 clAEAKO2_0#clCZWK1K_0#a_12_41# D GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#0 VCC clAEAKO2_0#clCZWK1K_0#Y clAEAKO2_0#clCZWK1K_1#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#1 clAEAKO2_0#clCZWK1K_1#a_18_54# clAEAKO2_0#clCZWK1K_1#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#2 clAEAKO2_0#Y clAEAKO2_0#clCZWK1K_1#a_2_6# clAEAKO2_0#clCZWK1K_1#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#3 clAEAKO2_0#clCZWK1K_1#a_35_54# clAEAKO2_0#clCZWK1K_0#Y clAEAKO2_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#4 VCC B clAEAKO2_0#clCZWK1K_1#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#5 clAEAKO2_0#clCZWK1K_1#a_12_41# B VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#6 GND clAEAKO2_0#clCZWK1K_0#Y clAEAKO2_0#clCZWK1K_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#7 clAEAKO2_0#clCZWK1K_1#a_18_6# clAEAKO2_0#clCZWK1K_1#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#8 clAEAKO2_0#Y clAEAKO2_0#clCZWK1K_0#Y clAEAKO2_0#clCZWK1K_1#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#9 clAEAKO2_0#clCZWK1K_1#a_35_6# clAEAKO2_0#clCZWK1K_1#a_2_6# clAEAKO2_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#10 GND B clAEAKO2_0#clCZWK1K_1#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_0#clCZWK1K_1#11 clAEAKO2_0#clCZWK1K_1#a_12_41# B GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_1#0 Y clAEAKO2_0#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_1#1 VCC A Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_1#2 clAEAKO2_1#a_9_6# clAEAKO2_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclAEAKO2_1#3 Y A clAEAKO2_1#a_9_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 3|4|NAND2X1|VOTER_G0_9_10=1|INPUT:Y-NAND2X1:A,B=1|INPUT:Y-VOTER_G0_9_10:A,B,C=3|VOTER_G0_9_10:Y-NAND2X1:A,B=1|111101
* 416 occurrences in design
* each contains 2 cells
* pin map: {'n6456': 'A', 'x721': 'B', 'x722': 'C', 'x723': 'D'} {'n6457': 'Y'}
* function: ~A|(B&C&~D)|(B&D&~C)|(C&D&~B)|(~B&~C&~D)
* Example occurence:
*   .subckt VOTER_G0_9_10 A=x721 B=x722 C=x723 Y=n6455
*   .subckt NAND2X1 A=n6455 B=n6456 Y=n6457
