.SUBCKT ROUTER_G4_30_104 A B Y VCC GND
MclPJDTIL_0#0 clPJDTIL_0#Y B VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPJDTIL_0#1 clPJDTIL_0#Y B GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPJDTIL_1#0 Y clPJDTIL_0#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPJDTIL_1#1 VCC A Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPJDTIL_1#2 clPJDTIL_1#a_9_6# clPJDTIL_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPJDTIL_1#3 Y A clPJDTIL_1#a_9_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 2|2|NAND2X1|INVX1=1|INPUT:Y-INVX1:A=1|INPUT:Y-NAND2X1:A,B=1|INVX1:Y-NAND2X1:A,B=1|1110
* 12 occurrences in design
* each contains 2 cells
* pin map: {'n66': 'A', 'x9': 'B'} {'n97': 'Y'}
* function: B|~A
* Example occurence:
*   .subckt INVX1 A=x9 Y=n65
*   .subckt NAND2X1 A=n65 B=n66 Y=n97
