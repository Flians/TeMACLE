.SUBCKT BAR_G0_0_1742 A B Y VCC GND
MclKERZGT_0#0 clKERZGT_0#Y B VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclKERZGT_0#1 clKERZGT_0#Y B GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclKERZGT_1#0 Y clKERZGT_0#Y VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclKERZGT_1#1 VCC A Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclKERZGT_1#2 clKERZGT_1#a_9_6# clKERZGT_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclKERZGT_1#3 Y A clKERZGT_1#a_9_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 2|2|NAND2X1|INVX1=1|INPUT:Y-INVX1:A=1|INPUT:Y-NAND2X1:A,B=1|INVX1:Y-NAND2X1:A,B=1|1110
* 120 occurrences in design
* each contains 2 cells
* pin map: {'n1506': 'A', 'x133': 'B'} {'n1889': 'Y'}
* function: B|~A
* Example occurence:
*   .subckt INVX1 A=x133 Y=n267
*   .subckt NAND2X1 A=n267 B=n1506 Y=n1889
