.SUBCKT ADDER_G2_0_605 A B C Y VCC GND
MclOFJ1YE_0#0 clOFJ1YE_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_0#1 clOFJ1YE_0#Y C GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#0 VCC B clOFJ1YE_1#cl7AM7QI_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#1 clOFJ1YE_1#cl7AM7QI_0#a_18_54# clOFJ1YE_1#cl7AM7QI_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#2 clOFJ1YE_1#cl7AM7QI_0#Y clOFJ1YE_1#cl7AM7QI_0#a_2_6# clOFJ1YE_1#cl7AM7QI_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#3 clOFJ1YE_1#cl7AM7QI_0#a_35_54# B clOFJ1YE_1#cl7AM7QI_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#4 VCC A clOFJ1YE_1#cl7AM7QI_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#5 clOFJ1YE_1#cl7AM7QI_0#a_12_41# A VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#6 GND B clOFJ1YE_1#cl7AM7QI_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#7 clOFJ1YE_1#cl7AM7QI_0#a_18_6# clOFJ1YE_1#cl7AM7QI_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#8 clOFJ1YE_1#cl7AM7QI_0#Y B clOFJ1YE_1#cl7AM7QI_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#9 clOFJ1YE_1#cl7AM7QI_0#a_35_6# clOFJ1YE_1#cl7AM7QI_0#a_2_6# clOFJ1YE_1#cl7AM7QI_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#10 GND A clOFJ1YE_1#cl7AM7QI_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_0#11 clOFJ1YE_1#cl7AM7QI_0#a_12_41# A GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#0 VCC clOFJ1YE_1#cl7AM7QI_0#Y clOFJ1YE_1#cl7AM7QI_1#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#1 clOFJ1YE_1#cl7AM7QI_1#a_18_54# clOFJ1YE_1#cl7AM7QI_1#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#2 Y clOFJ1YE_1#cl7AM7QI_1#a_2_6# clOFJ1YE_1#cl7AM7QI_1#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#3 clOFJ1YE_1#cl7AM7QI_1#a_35_54# clOFJ1YE_1#cl7AM7QI_0#Y Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#4 VCC clOFJ1YE_0#Y clOFJ1YE_1#cl7AM7QI_1#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#5 clOFJ1YE_1#cl7AM7QI_1#a_12_41# clOFJ1YE_0#Y VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#6 GND clOFJ1YE_1#cl7AM7QI_0#Y clOFJ1YE_1#cl7AM7QI_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#7 clOFJ1YE_1#cl7AM7QI_1#a_18_6# clOFJ1YE_1#cl7AM7QI_1#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#8 Y clOFJ1YE_1#cl7AM7QI_0#Y clOFJ1YE_1#cl7AM7QI_1#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#9 clOFJ1YE_1#cl7AM7QI_1#a_35_6# clOFJ1YE_1#cl7AM7QI_1#a_2_6# Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#10 GND clOFJ1YE_0#Y clOFJ1YE_1#cl7AM7QI_1#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclOFJ1YE_1#cl7AM7QI_1#11 clOFJ1YE_1#cl7AM7QI_1#a_12_41# clOFJ1YE_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 3|3|ADDER_G0_454_455|INVX1=1|INPUT:Y-ADDER_G0_454_455:A,B,C=2|INPUT:Y-INVX1:A=1|INVX1:Y-ADDER_G0_454_455:A,B,C=1|01111
* 33 occurrences in design
* each contains 2 cells
* pin map: {'x254': 'A', 'n732': 'B', 'x126': 'C'} {'y127': 'Y'}
* function: (A&B&~C)|(A&C&~B)|(B&C&~A)|(~A&~B&~C)
* Example occurence:
*   .subckt INVX1 A=x126 Y=n322
*   .subckt ADDER_G0_454_455 A=n322 B=x254 C=n732 Y=y127
