.SUBCKT ADDER_G2_0_605 A B C Y VCC GND
MclCK2XCA_0#0 clCK2XCA_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_0#1 clCK2XCA_0#Y C GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#0 VCC B clCK2XCA_1#clNF429V_0#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#1 clCK2XCA_1#clNF429V_0#a_18_54# clCK2XCA_1#clNF429V_0#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#2 clCK2XCA_1#clNF429V_0#Y clCK2XCA_1#clNF429V_0#a_2_6# clCK2XCA_1#clNF429V_0#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#3 clCK2XCA_1#clNF429V_0#a_35_54# B clCK2XCA_1#clNF429V_0#Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#4 VCC A clCK2XCA_1#clNF429V_0#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#5 clCK2XCA_1#clNF429V_0#a_12_41# A VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#6 GND B clCK2XCA_1#clNF429V_0#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#7 clCK2XCA_1#clNF429V_0#a_18_6# clCK2XCA_1#clNF429V_0#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#8 clCK2XCA_1#clNF429V_0#Y B clCK2XCA_1#clNF429V_0#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#9 clCK2XCA_1#clNF429V_0#a_35_6# clCK2XCA_1#clNF429V_0#a_2_6# clCK2XCA_1#clNF429V_0#Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#10 GND A clCK2XCA_1#clNF429V_0#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_0#11 clCK2XCA_1#clNF429V_0#a_12_41# A GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#0 VCC clCK2XCA_1#clNF429V_0#Y clCK2XCA_1#clNF429V_1#a_2_6# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#1 clCK2XCA_1#clNF429V_1#a_18_54# clCK2XCA_1#clNF429V_1#a_12_41# VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#2 Y clCK2XCA_1#clNF429V_1#a_2_6# clCK2XCA_1#clNF429V_1#a_18_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#3 clCK2XCA_1#clNF429V_1#a_35_54# clCK2XCA_1#clNF429V_0#Y Y VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#4 VCC clCK2XCA_0#Y clCK2XCA_1#clNF429V_1#a_35_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#5 clCK2XCA_1#clNF429V_1#a_12_41# clCK2XCA_0#Y VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#6 GND clCK2XCA_1#clNF429V_0#Y clCK2XCA_1#clNF429V_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#7 clCK2XCA_1#clNF429V_1#a_18_6# clCK2XCA_1#clNF429V_1#a_12_41# GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#8 Y clCK2XCA_1#clNF429V_0#Y clCK2XCA_1#clNF429V_1#a_18_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#9 clCK2XCA_1#clNF429V_1#a_35_6# clCK2XCA_1#clNF429V_1#a_2_6# Y GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#10 GND clCK2XCA_0#Y clCK2XCA_1#clNF429V_1#a_35_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclCK2XCA_1#clNF429V_1#11 clCK2XCA_1#clNF429V_1#a_12_41# clCK2XCA_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 3|3|ADDER_G0_454_455|INVX1=1|INPUT:Y-ADDER_G0_454_455:A,B,C=2|INPUT:Y-INVX1:A=1|INVX1:Y-ADDER_G0_454_455:A,B,C=1|01111
* 33 occurrences in design
* each contains 2 cells
* pin map: {'x254': 'A', 'n732': 'B', 'x126': 'C'} {'y127': 'Y'}
* function: (A&B&~C)|(A&C&~B)|(B&C&~A)|(~A&~B&~C)
* Example occurence:
*   .subckt INVX1 A=x126 Y=n322
*   .subckt ADDER_G0_454_455 A=n322 B=x254 C=n732 Y=y127
