.subckt COMPLEX25 cl4#vdd cl1#B cl2#B cl3#A cl5#Y cl4#gnd cl4#B cl3#gnd cl1#gnd cl5#vdd cl3#B cl0#vdd cl5#A cl1#A cl0#gnd cl2#A cl5#gnd cl1#vdd cl4#A cl2#vdd cl2#gnd cl3#vdd
Mcl0#0 cl0#Y cl1#Y cl0#vdd cl0#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0#1 cl0#vdd cl2#Y cl0#Y cl0#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0#2 cl0#Y cl3#Y cl0#vdd cl0#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0#3 cl0#a_9_6# cl1#Y cl0#gnd cl0#gnd nmos w=0.75u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0#4 cl0#a_14_6# cl2#Y cl0#a_9_6# cl0#gnd nmos w=0.75u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl0#5 cl0#Y cl3#Y cl0#a_14_6# cl0#gnd nmos w=0.75u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl1#0 cl1#Y cl1#A cl1#vdd cl1#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl1#1 cl1#vdd cl1#B cl1#Y cl1#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl1#2 cl1#a_9_6# cl1#A cl1#gnd cl1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl1#3 cl1#Y cl1#B cl1#a_9_6# cl1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl2#0 cl2#Y cl2#A cl2#vdd cl2#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl2#1 cl2#vdd cl2#B cl2#Y cl2#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl2#2 cl2#a_9_6# cl2#A cl2#gnd cl2#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl2#3 cl2#Y cl2#B cl2#a_9_6# cl2#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl3#0 cl3#Y cl3#A cl3#vdd cl3#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl3#1 cl3#vdd cl3#B cl3#Y cl3#vdd pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl3#2 cl3#a_9_6# cl3#A cl3#gnd cl3#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl3#3 cl3#Y cl3#B cl3#a_9_6# cl3#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl4#0 cl4#vdd cl4#A cl4#a_2_54# cl4#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl4#1 cl4#a_2_54# cl4#B cl4#vdd cl4#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl4#2 cl4#Y cl0#Y cl4#a_2_54# cl4#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl4#3 cl4#a_12_6# cl4#A cl4#gnd cl4#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl4#4 cl4#Y cl4#B cl4#a_12_6# cl4#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl4#5 cl4#gnd cl0#Y cl4#Y cl4#gnd nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#0 cl5#vdd cl5#A cl5#a_2_6# cl5#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#1 cl5#a_18_54# cl5#a_12_41# cl5#vdd cl5#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#2 cl5#Y cl5#a_2_6# cl5#a_18_54# cl5#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#3 cl5#a_35_54# cl5#A cl5#Y cl5#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#4 cl5#vdd cl4#Y cl5#a_35_54# cl5#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#5 cl5#a_12_41# cl4#Y cl5#vdd cl5#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#6 cl5#gnd cl5#A cl5#a_2_6# cl5#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#7 cl5#a_18_6# cl5#a_12_41# cl5#gnd cl5#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#8 cl5#Y cl5#A cl5#a_18_6# cl5#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#9 cl5#a_35_6# cl5#a_2_6# cl5#Y cl5#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#10 cl5#gnd cl4#Y cl5#a_35_6# cl5#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl5#11 cl5#a_12_41# cl4#Y cl5#gnd cl5#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ends COMPLEX25
* pattern code: [NAND3X1,NAND2X1,NAND2X1,NAND2X1]+AOI21X1_c0o0+XNOR2X1_c4o0
* 450 occurrences in design 
* each contains 6 cells
* Example occurence:
*   .subckt NAND3X1 A=n3887 B=n3888 C=n3889 Y=n3890
*   .subckt NAND2X1 A=n1464 B=n3416 Y=n3887
*   .subckt NAND2X1 A=n1372 B=n3471 Y=n3888
*   .subckt NAND2X1 A=n1295 B=n3765 Y=n3889
*   .subckt AOI21X1 A=n3423 B=n3592 C=n3890 Y=n3891
*   .subckt XNOR2X1 A=n63 B=n3891 Y=n3892
