.SUBCKT BAR_G3_1_2 A B C VDD VSS Y
MclJG59IU_0#M0 clJG59IU_0#Y C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_0#M1 clJG59IU_0#Y C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_1#clEHB6JD_0#M3 clJG59IU_1#clEHB6JD_0#net16 clJG59IU_0#Y VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MclJG59IU_1#clEHB6JD_0#M2 clJG59IU_1#clEHB6JD_0#Y A clJG59IU_1#clEHB6JD_0#net16 VSS nmos_lvt w=162.00n l=20n nfin=6
MclJG59IU_1#clEHB6JD_0#M1 clJG59IU_1#clEHB6JD_0#Y A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_1#clEHB6JD_0#M0 clJG59IU_1#clEHB6JD_0#Y clJG59IU_0#Y VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_1#clEHB6JD_1#cl0ODER2_0#M5 VSS clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net7 clJG59IU_1#clEHB6JD_1#cl0ODER2_0#Y VSS nmos_lvt w=162.00n l=20n nfin=6
MclJG59IU_1#clEHB6JD_1#cl0ODER2_0#M1 VSS clJG59IU_1#clEHB6JD_1#C clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MclJG59IU_1#clEHB6JD_1#cl0ODER2_0#M2 VSS B clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MclJG59IU_1#clEHB6JD_1#cl0ODER2_0#M0 VDD clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net7 clJG59IU_1#clEHB6JD_1#cl0ODER2_0#Y VDD pmos_lvt w=162.00n l=20n nfin=6
MclJG59IU_1#clEHB6JD_1#cl0ODER2_0#M4 clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net15 clJG59IU_1#clEHB6JD_1#C clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net7 VDD pmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_1#clEHB6JD_1#cl0ODER2_0#M3 VDD B clJG59IU_1#clEHB6JD_1#cl0ODER2_0#net15 VDD pmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_1#clEHB6JD_1#cl0ODER2_1#M4 Y clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net10 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MclJG59IU_1#clEHB6JD_1#cl0ODER2_1#M1 clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net10 clJG59IU_1#clEHB6JD_0#Y VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MclJG59IU_1#clEHB6JD_1#cl0ODER2_1#M0 clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net10 clJG59IU_1#clEHB6JD_1#cl0ODER2_0#Y VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MclJG59IU_1#clEHB6JD_1#cl0ODER2_1#M5 Y clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net10 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MclJG59IU_1#clEHB6JD_1#cl0ODER2_1#M3 clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net20 clJG59IU_1#clEHB6JD_1#cl0ODER2_0#Y VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MclJG59IU_1#clEHB6JD_1#cl0ODER2_1#M2 clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net10 clJG59IU_1#clEHB6JD_0#Y clJG59IU_1#clEHB6JD_1#cl0ODER2_1#net20 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS 
* pattern code: 4|3|BAR_G2_3_5|INVx1=1|INPUT:Y-BAR_G2_3_5:A=1|INPUT:Y-BAR_G2_3_5:B=1|INPUT:Y-INVx1:A=1|INVx1:Y-BAR_G2_3_5:C=1|01111
* 65 occurrences in design
* each contains 2 cells
* function: (A&C)|(B&~A)
* Example occurence:
*   .subckt INVx1 A=x58 Y=n188
*   .subckt BAR_G2_3_5 A=x57 B=n250 C=n188 Y=n358
