.SUBCKT CAVLC_G4_0_152 A B C Y VCC GND
Mcl6DO165_0#0 cl6DO165_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_0#1 cl6DO165_0#Y C GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_1#0 VCC cl6DO165_0#Y cl6DO165_1#a_2_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_1#1 cl6DO165_1#a_2_54# A VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_1#2 Y B cl6DO165_1#a_2_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_1#3 cl6DO165_1#a_12_6# cl6DO165_0#Y GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_1#4 Y A cl6DO165_1#a_12_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
Mcl6DO165_1#5 GND B Y GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 2|3|AOI21X1|INVX1=1|INPUT:Y-AOI21X1:A,B=1|INPUT:Y-AOI21X1:C=1|INPUT:Y-INVX1:A=1|INVX1:Y-AOI21X1:A,B=1|01111
* 28 occurrences in design
* each contains 2 cells
* pin map: {'n158': 'A', 'n154': 'B', 'x0': 'C'} {'n159': 'Y'}
* function: ~B&(C|~A)
* Example occurence:
*   .subckt INVX1 A=x0 Y=n12
*   .subckt AOI21X1 A=n12 B=n158 C=n154 Y=n159
