.SUBCKT SQRT_G0_173_198_231 A B C Y VCC GND
MclPVOFZ6_0#0 clPVOFZ6_0#vdd C clPVOFZ6_0#a_2_6# clPVOFZ6_0#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#1 clPVOFZ6_0#a_18_54# clPVOFZ6_0#a_12_41# clPVOFZ6_0#vdd clPVOFZ6_0#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#2 clPVOFZ6_0#Y clPVOFZ6_0#a_2_6# clPVOFZ6_0#a_18_54# clPVOFZ6_0#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#3 clPVOFZ6_0#a_35_54# C clPVOFZ6_0#Y clPVOFZ6_0#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#4 clPVOFZ6_0#vdd B clPVOFZ6_0#a_35_54# clPVOFZ6_0#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#5 clPVOFZ6_0#a_12_41# B clPVOFZ6_0#vdd clPVOFZ6_0#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#6 clPVOFZ6_0#gnd C clPVOFZ6_0#a_2_6# clPVOFZ6_0#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#7 clPVOFZ6_0#a_18_6# clPVOFZ6_0#a_12_41# clPVOFZ6_0#gnd clPVOFZ6_0#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#8 clPVOFZ6_0#Y C clPVOFZ6_0#a_18_6# clPVOFZ6_0#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#9 clPVOFZ6_0#a_35_6# clPVOFZ6_0#a_2_6# clPVOFZ6_0#Y clPVOFZ6_0#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#10 clPVOFZ6_0#gnd B clPVOFZ6_0#a_35_6# clPVOFZ6_0#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_0#11 clPVOFZ6_0#a_12_41# B clPVOFZ6_0#gnd clPVOFZ6_0#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#0 clPVOFZ6_1#vdd clPVOFZ6_0#Y clPVOFZ6_1#a_2_6# clPVOFZ6_1#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#1 clPVOFZ6_1#a_18_54# clPVOFZ6_1#a_13_43# clPVOFZ6_1#vdd clPVOFZ6_1#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#2 Y clPVOFZ6_0#Y clPVOFZ6_1#a_18_54# clPVOFZ6_1#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#3 clPVOFZ6_1#a_35_54# clPVOFZ6_1#a_2_6# Y clPVOFZ6_1#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#4 clPVOFZ6_1#vdd A clPVOFZ6_1#a_35_54# clPVOFZ6_1#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#5 clPVOFZ6_1#a_13_43# A clPVOFZ6_1#vdd clPVOFZ6_1#vdd pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#6 clPVOFZ6_1#gnd clPVOFZ6_0#Y clPVOFZ6_1#a_2_6# clPVOFZ6_1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#7 clPVOFZ6_1#a_18_6# clPVOFZ6_1#a_13_43# clPVOFZ6_1#gnd clPVOFZ6_1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#8 Y clPVOFZ6_1#a_2_6# clPVOFZ6_1#a_18_6# clPVOFZ6_1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#9 clPVOFZ6_1#a_35_6# clPVOFZ6_0#Y Y clPVOFZ6_1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#10 clPVOFZ6_1#gnd A clPVOFZ6_1#a_35_6# clPVOFZ6_1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclPVOFZ6_1#11 clPVOFZ6_1#a_13_43# A clPVOFZ6_1#gnd clPVOFZ6_1#gnd nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS
* pattern code: 3|3|XNOR2X1|INVX1=1|XNOR2X1=1|INPUT:Y-XNOR2X1:A,B=3|INVX1:Y-XNOR2X1:A,B=1|XNOR2X1:Y-INVX1:A=1|111101
* 1493 occurrences in design
* each contains 3 cells
* pin map: {'n488': 'A', 'n417': 'B', 'n350': 'C'} {'n489': 'Y'}
* function: (A&B&~C)|(A&C&~B)|(B&C&~A)|(~A&~B&~C)
* Example occurence:
*   .subckt XNOR2X1 A=n417 B=n350 Y=n418
*   .subckt INVX1 A=n418 Y=n419
*   .subckt XNOR2X1 A=n488 B=n419 Y=n489
