.SUBCKT SQUARE_G2_2_28 A B C Y VCC GND
MclWA32Y5_0#0 clWA32Y5_0#Y C VCC VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_0#1 clWA32Y5_0#Y C GND GND nmos w=0.25u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_1#0 clWA32Y5_1#a_9_54# clWA32Y5_0#Y VCC VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_1#1 Y A clWA32Y5_1#a_9_54# VCC pmos w=1u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_1#2 VCC B Y VCC pmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_1#3 GND clWA32Y5_0#Y clWA32Y5_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_1#4 clWA32Y5_1#a_2_6# A GND GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
MclWA32Y5_1#5 Y B clWA32Y5_1#a_2_6# GND nmos w=0.5u l=0.05u
+ ad=0p pd=0u as=0p ps=0u
.ENDS 
* pattern code: 2|3|OAI21X1|INVX1=1|INPUT:Y-INVX1:A=1|INPUT:Y-OAI21X1:A,B=1|INPUT:Y-OAI21X1:C=1|INVX1:Y-OAI21X1:A,B=1|11110
* 921 occurrences in design
* each contains 2 cells
* pin map: {'n70': 'A', 'n152': 'B', 'x1': 'C'} {'n153': 'Y'}
* function: ~B|(C&~A)
* Example occurence:
*   .subckt INVX1 A=x1 Y=n67
*   .subckt OAI21X1 A=n67 B=n70 C=n152 Y=n153
